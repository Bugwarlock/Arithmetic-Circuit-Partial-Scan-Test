
//Verilog file of module fourFunc


`timescale 1 ns / 1ns

module fourFunc_net_Unfolded(clk,
rst,
start,
func,
x,
//ppIn
PPI0 ,
PPI1 ,
PPI2 ,
PPI3 ,
PPI4 ,
PPI5 ,
PPI6 ,
PPI7 ,
PPI8 ,
PPI9 ,
PPI10,
PPI11,
PPI12,
PPI13,
PPI14,
PPI15,
PPI16,
PPI17,
PPI18,
PPI19,
PPI20,
PPI21,
PPI22,
PPI23,
PPI24,
PPI25,
PPI26,
PPI27,
PPI28,
PPI29,
PPI30,
PPI31,
PPI32,
PPI33,
PPI34,
PPI35,
PPI36,
//ppIn
busy,
resultIPart,
resultFPart,
//ppOut

PPO0 ,
PPO1 ,
PPO2 ,
PPO3 ,
PPO4 ,
PPO5 ,
PPO6 ,
PPO7 ,
PPO8 ,
PPO9 ,
PPO10,
PPO11,
PPO12,
PPO13,
PPO14,
PPO15,
PPO16,
PPO17,
PPO18,
PPO19,
PPO20,
PPO21,
PPO22,
PPO23,
PPO24,
PPO25,
PPO26,
PPO27,
PPO28,
PPO29,
PPO30,
PPO31,
PPO32,
PPO33,
PPO34,
PPO35,
PPO36);


	input	clk;
	input	rst;
	input	start;
input [0:1]func;
input [0:7]x;
/////
input PPI0 ;
input PPI1 ;
input PPI2 ;
input PPI3 ;
input PPI4 ;
input PPI5 ;
input PPI6 ;
input PPI7 ;
input PPI8 ;
input PPI9 ;
input PPI10;
input PPI11;
input PPI12;
input PPI13;
input PPI14;
input PPI15;
input PPI16;
input PPI17;
input PPI18;
input PPI19;
input PPI20;
input PPI21;
input PPI22;
input PPI23;
input PPI24;
input PPI25;
input PPI26;
input PPI27;
input PPI28;
input PPI29;
input PPI30;
input PPI31;
input PPI32;
input PPI33;
input PPI34;
input PPI35;
input PPI36;
////
	output 	busy;
output [0:1]resultIPart;
output [0:7]resultFPart;
//// 
output PPO0 ;
output PPO1 ;
output PPO2 ;
output PPO3 ;
output PPO4 ;
output PPO5 ;
output PPO6 ;
output PPO7 ;
output PPO8 ;
output PPO9 ;
output PPO10;
output PPO11;
output PPO12;
output PPO13;
output PPO14;
output PPO15;
output PPO16;
output PPO17;
output PPO18;
output PPO19;
output PPO20;
output PPO21;
output PPO22;
output PPO23;
output PPO24;
output PPO25;
output PPO26;
output PPO27;
output PPO28;
output PPO29;
output PPO30;
output PPO31;
output PPO32;
output PPO33;
output PPO34;
output PPO35;
output PPO36;
///
wire
fourFunc_wire_1,
fourFunc_wire_2,
fourFunc_wire_3,
fourFunc_wire_4,
fourFunc_wire_5,
fourFunc_wire_6,
fourFunc_wire_7,
fourFunc_wire_8,
fourFunc_wire_9,
fourFunc_wire_10,
fourFunc_wire_11,
fourFunc_wire_12,
fourFunc_wire_13,
fourFunc_wire_14,
fourFunc_wire_15,
fourFunc_wire_16,
fourFunc_wire_17,
fourFunc_wire_18,
fourFunc_wire_19,
fourFunc_wire_20,
fourFunc_wire_21,
fourFunc_wire_22,
fourFunc_wire_23,
fourFunc_wire_24,
fourFunc_wire_25,
fourFunc_wire_26,
fourFunc_wire_27,
fourFunc_wire_28,
fourFunc_wire_29,
fourFunc_wire_30,
fourFunc_wire_31,
fourFunc_wire_32,
fourFunc_wire_33,
fourFunc_wire_34,
fourFunc_wire_35,
fourFunc_wire_36,
fourFunc_wire_37,
fourFunc_wire_38,
fourFunc_wire_39,
fourFunc_wire_40,
fourFunc_wire_41,
fourFunc_wire_42,
fourFunc_wire_43,
fourFunc_wire_44,
fourFunc_wire_45,
fourFunc_wire_46,
fourFunc_wire_47,
fourFunc_wire_48,
fourFunc_wire_49,
fourFunc_wire_50,
fourFunc_wire_51,
fourFunc_wire_52,
fourFunc_wire_53,
fourFunc_wire_54,
fourFunc_wire_55,
fourFunc_wire_56,
fourFunc_wire_57,
fourFunc_wire_58,
fourFunc_wire_59,
fourFunc_wire_60,
fourFunc_wire_61,
fourFunc_wire_62,
fourFunc_wire_63,
fourFunc_wire_64,
fourFunc_wire_65,
fourFunc_wire_66,
fourFunc_wire_67,
fourFunc_wire_68,
fourFunc_wire_69,
fourFunc_wire_70,
fourFunc_wire_71,
fourFunc_wire_72,
fourFunc_wire_73,
fourFunc_wire_74,
fourFunc_wire_75,
fourFunc_wire_76,
fourFunc_wire_77,
fourFunc_wire_78,
fourFunc_wire_79,
fourFunc_wire_80,
fourFunc_wire_81,
fourFunc_wire_82,
fourFunc_wire_83,
fourFunc_wire_84,
fourFunc_wire_85,
fourFunc_wire_86,
fourFunc_wire_87,
fourFunc_wire_88,
fourFunc_wire_89,
fourFunc_wire_90,
fourFunc_wire_91,
fourFunc_wire_92,
fourFunc_wire_93,
fourFunc_wire_94,
fourFunc_wire_95,
fourFunc_wire_96,
fourFunc_wire_97,
fourFunc_wire_98,
fourFunc_wire_99,
fourFunc_wire_100,
fourFunc_wire_101,
fourFunc_wire_102,
fourFunc_wire_103,
fourFunc_wire_104,
fourFunc_wire_105,
fourFunc_wire_106,
fourFunc_wire_107,
fourFunc_wire_108,
fourFunc_wire_109,
fourFunc_wire_110,
fourFunc_wire_111,
fourFunc_wire_112,
fourFunc_wire_113,
fourFunc_wire_114,
fourFunc_wire_115,
fourFunc_wire_116,
fourFunc_wire_117,
fourFunc_wire_118,
fourFunc_wire_119,
fourFunc_wire_120,
fourFunc_wire_121,
fourFunc_wire_122,
fourFunc_wire_123,
fourFunc_wire_124,
fourFunc_wire_125,
fourFunc_wire_126,
fourFunc_wire_127,
fourFunc_wire_128,
fourFunc_wire_129,
fourFunc_wire_130,
fourFunc_wire_131,
fourFunc_wire_132,
fourFunc_wire_133,
fourFunc_wire_134,
fourFunc_wire_135,
fourFunc_wire_136,
fourFunc_wire_137,
fourFunc_wire_138,
fourFunc_wire_139,
fourFunc_wire_140,
fourFunc_wire_141,
fourFunc_wire_142,
fourFunc_wire_143,
fourFunc_wire_144,
fourFunc_wire_145,
fourFunc_wire_146,
fourFunc_wire_147,
fourFunc_wire_148,
fourFunc_wire_149,
fourFunc_wire_150,
fourFunc_wire_151,
fourFunc_wire_152,
fourFunc_wire_153,
fourFunc_wire_154,
fourFunc_wire_155,
fourFunc_wire_156,
fourFunc_wire_157,
fourFunc_wire_158,
fourFunc_wire_159,
fourFunc_wire_160,
fourFunc_wire_161,
fourFunc_wire_162,
fourFunc_wire_163,
fourFunc_wire_164,
fourFunc_wire_165,
fourFunc_wire_166,
fourFunc_wire_167,
fourFunc_wire_168,
fourFunc_wire_169,
fourFunc_wire_170,
fourFunc_wire_171,
fourFunc_wire_172,
fourFunc_wire_173,
fourFunc_wire_174,
fourFunc_wire_175,
fourFunc_wire_176,
fourFunc_wire_177,
fourFunc_wire_178,
fourFunc_wire_179,
fourFunc_wire_180,
fourFunc_wire_181,
fourFunc_wire_182,
fourFunc_wire_183,
fourFunc_wire_184,
fourFunc_wire_185,
fourFunc_wire_186,
fourFunc_wire_187,
fourFunc_wire_188,
fourFunc_wire_189,
fourFunc_wire_190,
fourFunc_wire_191,
fourFunc_wire_192,
fourFunc_wire_193,
fourFunc_wire_194,
fourFunc_wire_195,
fourFunc_wire_196,
fourFunc_wire_197,
fourFunc_wire_198,
fourFunc_wire_199,
fourFunc_wire_200,
fourFunc_wire_201,
fourFunc_wire_202,
fourFunc_wire_203,
fourFunc_wire_204,
fourFunc_wire_205,
fourFunc_wire_206,
fourFunc_wire_207,
fourFunc_wire_208,
fourFunc_wire_209,
fourFunc_wire_210,
fourFunc_wire_211,
fourFunc_wire_212,
fourFunc_wire_213,
fourFunc_wire_214,
fourFunc_wire_215,
fourFunc_wire_216,
fourFunc_wire_217,
fourFunc_wire_218,
fourFunc_wire_219,
fourFunc_wire_220,
fourFunc_wire_221,
fourFunc_wire_222,
fourFunc_wire_223,
fourFunc_wire_224,
fourFunc_wire_225,
fourFunc_wire_226,
fourFunc_wire_227,
fourFunc_wire_228,
fourFunc_wire_229,
fourFunc_wire_230,
fourFunc_wire_231,
fourFunc_wire_232,
fourFunc_wire_233,
fourFunc_wire_234,
fourFunc_wire_235,
fourFunc_wire_236,
fourFunc_wire_237,
fourFunc_wire_238,
fourFunc_wire_239,
fourFunc_wire_240,
fourFunc_wire_241,
fourFunc_wire_242,
fourFunc_wire_243,
fourFunc_wire_244,
fourFunc_wire_245,
fourFunc_wire_246,
fourFunc_wire_247,
fourFunc_wire_248,
fourFunc_wire_249,
fourFunc_wire_250,
fourFunc_wire_251,
fourFunc_wire_252,
fourFunc_wire_253,
fourFunc_wire_254,
fourFunc_wire_255,
fourFunc_wire_256,
fourFunc_wire_257,
fourFunc_wire_258,
fourFunc_wire_259,
fourFunc_wire_260,
fourFunc_wire_261,
fourFunc_wire_262,
fourFunc_wire_263,
fourFunc_wire_264,
fourFunc_wire_265,
fourFunc_wire_266,
fourFunc_wire_267,
fourFunc_wire_268,
fourFunc_wire_269,
fourFunc_wire_270,
fourFunc_wire_271,
fourFunc_wire_272,
fourFunc_wire_273,
fourFunc_wire_274,
fourFunc_wire_275,
fourFunc_wire_276,
fourFunc_wire_277,
fourFunc_wire_278,
fourFunc_wire_279,
fourFunc_wire_280,
fourFunc_wire_281,
fourFunc_wire_282,
fourFunc_wire_283,
fourFunc_wire_284,
fourFunc_wire_285,
fourFunc_wire_286,
fourFunc_wire_287,
fourFunc_wire_288,
fourFunc_wire_289,
fourFunc_wire_290,
fourFunc_wire_291,
fourFunc_wire_292,
fourFunc_wire_293,
fourFunc_wire_294,
fourFunc_wire_295,
fourFunc_wire_296,
fourFunc_wire_297,
fourFunc_wire_298,
fourFunc_wire_299,
fourFunc_wire_300,
fourFunc_wire_301,
fourFunc_wire_302,
fourFunc_wire_303,
fourFunc_wire_304,
fourFunc_wire_305,
fourFunc_wire_306,
fourFunc_wire_307,
fourFunc_wire_308,
fourFunc_wire_309,
fourFunc_wire_310,
fourFunc_wire_311,
fourFunc_wire_312,
fourFunc_wire_313,
fourFunc_wire_314,
fourFunc_wire_315,
fourFunc_wire_316,
fourFunc_wire_317,
fourFunc_wire_318,
fourFunc_wire_319,
fourFunc_wire_320,
fourFunc_wire_321,
fourFunc_wire_322,
fourFunc_wire_323,
fourFunc_wire_324,
fourFunc_wire_325,
fourFunc_wire_326,
fourFunc_wire_327,
fourFunc_wire_328,
fourFunc_wire_329,
fourFunc_wire_330,
fourFunc_wire_331,
fourFunc_wire_332,
fourFunc_wire_333,
fourFunc_wire_334,
fourFunc_wire_335,
fourFunc_wire_336,
fourFunc_wire_337,
fourFunc_wire_338,
fourFunc_wire_339,
fourFunc_wire_340,
fourFunc_wire_341,
fourFunc_wire_342,
fourFunc_wire_343,
fourFunc_wire_344,
fourFunc_wire_345,
fourFunc_wire_346,
fourFunc_wire_347,
fourFunc_wire_348,
fourFunc_wire_349,
fourFunc_wire_350,
fourFunc_wire_351,
fourFunc_wire_352,
fourFunc_wire_353,
fourFunc_wire_354,
fourFunc_wire_355,
fourFunc_wire_356,
fourFunc_wire_357,
fourFunc_wire_358,
fourFunc_wire_359,
fourFunc_wire_360,
fourFunc_wire_361,
fourFunc_wire_362,
fourFunc_wire_363,
fourFunc_wire_364,
fourFunc_wire_365,
fourFunc_wire_366,
fourFunc_wire_367,
fourFunc_wire_368,
fourFunc_wire_369,
fourFunc_wire_370,
fourFunc_wire_371,
fourFunc_wire_372,
fourFunc_wire_373,
fourFunc_wire_374,
fourFunc_wire_375,
fourFunc_wire_376,
fourFunc_wire_377,
fourFunc_wire_378,
fourFunc_wire_379,
fourFunc_wire_380,
fourFunc_wire_381,
fourFunc_wire_382,
fourFunc_wire_383,
fourFunc_wire_384,
fourFunc_wire_385,
fourFunc_wire_386,
fourFunc_wire_387,
fourFunc_wire_388,
fourFunc_wire_389,
fourFunc_wire_390,
fourFunc_wire_391,
fourFunc_wire_392,
fourFunc_wire_393,
fourFunc_wire_394,
fourFunc_wire_395,
fourFunc_wire_396,
fourFunc_wire_397,
fourFunc_wire_398,
fourFunc_wire_399,
fourFunc_wire_400,
fourFunc_wire_401,
fourFunc_wire_402,
fourFunc_wire_403,
fourFunc_wire_404,
fourFunc_wire_405,
fourFunc_wire_406,
fourFunc_wire_407,
fourFunc_wire_408,
fourFunc_wire_409,
fourFunc_wire_410,
fourFunc_wire_411,
fourFunc_wire_412,
fourFunc_wire_413,
fourFunc_wire_414,
fourFunc_wire_415,
fourFunc_wire_416,
fourFunc_wire_417,
fourFunc_wire_418,
fourFunc_wire_419,
fourFunc_wire_420,
fourFunc_wire_421,
fourFunc_wire_422,
fourFunc_wire_423,
fourFunc_wire_424,
fourFunc_wire_425,
fourFunc_wire_426,
fourFunc_wire_427,
fourFunc_wire_428,
fourFunc_wire_429,
fourFunc_wire_430,
fourFunc_wire_431,
fourFunc_wire_432,
fourFunc_wire_433,
fourFunc_wire_434,
fourFunc_wire_435,
fourFunc_wire_436,
fourFunc_wire_437,
fourFunc_wire_438,
fourFunc_wire_439,
fourFunc_wire_440,
fourFunc_wire_441,
fourFunc_wire_442,
fourFunc_wire_443,
fourFunc_wire_444,
fourFunc_wire_445,
fourFunc_wire_446,
fourFunc_wire_447,
fourFunc_wire_448,
fourFunc_wire_449,
fourFunc_wire_450,
fourFunc_wire_451,
fourFunc_wire_452,
fourFunc_wire_453,
fourFunc_wire_454,
fourFunc_wire_455,
fourFunc_wire_456,
fourFunc_wire_457,
fourFunc_wire_458,
fourFunc_wire_459,
fourFunc_wire_460,
fourFunc_wire_461,
fourFunc_wire_462,
fourFunc_wire_463,
fourFunc_wire_464,
fourFunc_wire_465,
fourFunc_wire_466,
fourFunc_wire_467,
fourFunc_wire_468,
fourFunc_wire_469,
fourFunc_wire_470,
fourFunc_wire_471,
fourFunc_wire_472,
fourFunc_wire_473,
fourFunc_wire_474,
fourFunc_wire_475,
fourFunc_wire_476,
fourFunc_wire_477,
fourFunc_wire_478,
fourFunc_wire_479,
fourFunc_wire_480,
fourFunc_wire_481,
fourFunc_wire_482,
fourFunc_wire_483,
fourFunc_wire_484,
fourFunc_wire_485,
fourFunc_wire_486,
fourFunc_wire_487,
fourFunc_wire_488,
fourFunc_wire_489,
fourFunc_wire_490,
fourFunc_wire_491,
fourFunc_wire_492,
fourFunc_wire_493,
fourFunc_wire_494,
fourFunc_wire_495,
fourFunc_wire_496,
fourFunc_wire_497,
fourFunc_wire_498,
fourFunc_wire_499,
fourFunc_wire_500,
fourFunc_wire_501,
fourFunc_wire_502,
fourFunc_wire_503,
fourFunc_wire_504,
fourFunc_wire_505,
fourFunc_wire_506,
fourFunc_wire_507,
fourFunc_wire_508,
fourFunc_wire_509,
fourFunc_wire_510,
fourFunc_wire_511,
fourFunc_wire_512,
fourFunc_wire_513,
fourFunc_wire_514,
fourFunc_wire_515,
fourFunc_wire_516,
fourFunc_wire_517,
fourFunc_wire_518,
fourFunc_wire_519,
fourFunc_wire_520,
fourFunc_wire_521,
fourFunc_wire_522,
fourFunc_wire_523,
fourFunc_wire_524,
fourFunc_wire_525,
fourFunc_wire_526,
fourFunc_wire_527,
fourFunc_wire_528,
fourFunc_wire_529,
fourFunc_wire_530,
fourFunc_wire_531,
fourFunc_wire_532,
fourFunc_wire_533,
fourFunc_wire_534,
fourFunc_wire_535,
fourFunc_wire_536,
fourFunc_wire_537,
fourFunc_wire_538,
fourFunc_wire_539,
fourFunc_wire_540,
fourFunc_wire_541,
fourFunc_wire_542,
fourFunc_wire_543,
fourFunc_wire_544,
fourFunc_wire_545,
fourFunc_wire_546,
fourFunc_wire_547,
fourFunc_wire_548,
fourFunc_wire_549,
fourFunc_wire_550,
fourFunc_wire_551,
fourFunc_wire_552,
fourFunc_wire_553,
fourFunc_wire_554,
fourFunc_wire_555,
fourFunc_wire_556,
fourFunc_wire_557,
fourFunc_wire_558,
fourFunc_wire_559,
fourFunc_wire_560,
fourFunc_wire_561,
fourFunc_wire_562,
fourFunc_wire_563,
fourFunc_wire_564,
fourFunc_wire_565,
fourFunc_wire_566,
fourFunc_wire_567,
fourFunc_wire_568,
fourFunc_wire_569,
fourFunc_wire_570,
fourFunc_wire_571,
fourFunc_wire_572,
fourFunc_wire_573,
fourFunc_wire_574,
fourFunc_wire_575,
fourFunc_wire_576,
fourFunc_wire_577,
fourFunc_wire_578,
fourFunc_wire_579,
fourFunc_wire_580,
fourFunc_wire_581,
fourFunc_wire_582,
fourFunc_wire_583,
fourFunc_wire_584,
fourFunc_wire_585,
fourFunc_wire_586,
fourFunc_wire_587,
fourFunc_wire_588,
fourFunc_wire_589,
fourFunc_wire_590,
fourFunc_wire_591,
fourFunc_wire_592,
fourFunc_wire_593,
fourFunc_wire_594,
fourFunc_wire_595,
fourFunc_wire_596,
fourFunc_wire_597,
fourFunc_wire_598,
fourFunc_wire_599,
fourFunc_wire_600,
fourFunc_wire_601,
fourFunc_wire_602,
fourFunc_wire_603,
fourFunc_wire_604,
fourFunc_wire_605,
fourFunc_wire_606,
fourFunc_wire_607,
fourFunc_wire_608,
fourFunc_wire_609,
fourFunc_wire_610,
fourFunc_wire_611,
fourFunc_wire_612,
fourFunc_wire_613,
fourFunc_wire_614,
fourFunc_wire_615,
fourFunc_wire_616,
fourFunc_wire_617,
fourFunc_wire_618,
fourFunc_wire_619,
fourFunc_wire_620,
fourFunc_wire_621,
fourFunc_wire_622,
fourFunc_wire_623,
fourFunc_wire_624,
fourFunc_wire_625,
fourFunc_wire_626,
fourFunc_wire_627,
fourFunc_wire_628,
fourFunc_wire_629,
fourFunc_wire_630,
fourFunc_wire_631,
fourFunc_wire_632,
fourFunc_wire_633,
fourFunc_wire_634,
fourFunc_wire_635,
fourFunc_wire_636,
fourFunc_wire_637,
fourFunc_wire_638,
fourFunc_wire_639,
fourFunc_wire_640,
fourFunc_wire_641,
fourFunc_wire_642,
fourFunc_wire_643,
fourFunc_wire_644,
fourFunc_wire_645,
fourFunc_wire_646,
fourFunc_wire_647,
fourFunc_wire_648,
fourFunc_wire_649,
fourFunc_wire_650,
fourFunc_wire_651,
fourFunc_wire_652,
fourFunc_wire_653,
fourFunc_wire_654,
fourFunc_wire_655,
fourFunc_wire_656,
fourFunc_wire_657,
fourFunc_wire_658,
fourFunc_wire_659,
fourFunc_wire_660,
fourFunc_wire_661,
fourFunc_wire_662,
fourFunc_wire_663,
fourFunc_wire_664,
fourFunc_wire_665,
fourFunc_wire_666,
fourFunc_wire_667,
fourFunc_wire_668,
fourFunc_wire_669,
fourFunc_wire_670,
fourFunc_wire_671,
fourFunc_wire_672,
fourFunc_wire_673,
fourFunc_wire_674,
fourFunc_wire_675,
fourFunc_wire_676,
fourFunc_wire_677,
fourFunc_wire_678,
fourFunc_wire_679,
fourFunc_wire_680,
fourFunc_wire_681,
fourFunc_wire_682,
fourFunc_wire_683,
fourFunc_wire_684,
fourFunc_wire_685,
fourFunc_wire_686,
fourFunc_wire_687,
fourFunc_wire_688,
fourFunc_wire_689,
fourFunc_wire_690,
fourFunc_wire_691,
fourFunc_wire_692,
fourFunc_wire_693,
fourFunc_wire_694,
fourFunc_wire_695,
fourFunc_wire_696,
fourFunc_wire_697,
fourFunc_wire_698,
fourFunc_wire_699,
fourFunc_wire_700,
fourFunc_wire_701,
fourFunc_wire_702,
fourFunc_wire_703,
fourFunc_wire_704,
fourFunc_wire_705,
fourFunc_wire_706,
fourFunc_wire_707,
fourFunc_wire_708,
fourFunc_wire_709,
fourFunc_wire_710,
fourFunc_wire_711,
fourFunc_wire_712,
fourFunc_wire_713,
fourFunc_wire_714,
fourFunc_wire_715,
fourFunc_wire_716,
fourFunc_wire_717,
fourFunc_wire_718,
fourFunc_wire_719,
fourFunc_wire_720,
fourFunc_wire_721,
fourFunc_wire_722,
fourFunc_wire_723,
fourFunc_wire_724,
fourFunc_wire_725,
fourFunc_wire_726,
fourFunc_wire_727,
fourFunc_wire_728,
fourFunc_wire_729,
fourFunc_wire_730,
fourFunc_wire_731,
fourFunc_wire_732,
fourFunc_wire_733,
fourFunc_wire_734,
fourFunc_wire_735,
fourFunc_wire_736,
fourFunc_wire_737,
fourFunc_wire_738,
fourFunc_wire_739,
fourFunc_wire_740,
fourFunc_wire_741,
fourFunc_wire_742,
fourFunc_wire_743,
fourFunc_wire_744,
fourFunc_wire_745,
fourFunc_wire_746,
fourFunc_wire_747,
fourFunc_wire_748,
fourFunc_wire_749,
fourFunc_wire_750,
fourFunc_wire_751,
fourFunc_wire_752,
fourFunc_wire_753,
fourFunc_wire_754,
fourFunc_wire_755,
fourFunc_wire_756,
fourFunc_wire_757,
fourFunc_wire_758,
fourFunc_wire_759,
fourFunc_wire_760,
fourFunc_wire_761,
fourFunc_wire_762,
fourFunc_wire_763,
fourFunc_wire_764,
fourFunc_wire_765,
fourFunc_wire_766,
fourFunc_wire_767,
fourFunc_wire_768,
fourFunc_wire_769,
fourFunc_wire_770,
fourFunc_wire_771,
fourFunc_wire_772,
fourFunc_wire_773,
fourFunc_wire_774,
fourFunc_wire_775,
fourFunc_wire_776,
fourFunc_wire_777,
fourFunc_wire_778,
fourFunc_wire_779,
fourFunc_wire_780,
fourFunc_wire_781,
fourFunc_wire_782,
fourFunc_wire_783,
fourFunc_wire_784,
fourFunc_wire_785,
fourFunc_wire_786,
fourFunc_wire_787,
fourFunc_wire_788,
fourFunc_wire_789,
fourFunc_wire_790,
fourFunc_wire_791,
fourFunc_wire_792,
fourFunc_wire_793,
fourFunc_wire_794,
fourFunc_wire_795,
fourFunc_wire_796,
fourFunc_wire_797,
fourFunc_wire_798,
fourFunc_wire_799,
fourFunc_wire_800,
fourFunc_wire_801,
fourFunc_wire_802,
fourFunc_wire_803,
fourFunc_wire_804,
fourFunc_wire_805,
fourFunc_wire_806,
fourFunc_wire_807,
fourFunc_wire_808,
fourFunc_wire_809,
fourFunc_wire_810,
fourFunc_wire_811,
fourFunc_wire_812,
fourFunc_wire_813,
fourFunc_wire_814,
fourFunc_wire_815,
fourFunc_wire_816,
fourFunc_wire_817,
fourFunc_wire_818,
fourFunc_wire_819,
fourFunc_wire_820,
fourFunc_wire_821,
fourFunc_wire_822,
fourFunc_wire_823,
fourFunc_wire_824,
fourFunc_wire_825,
fourFunc_wire_826,
fourFunc_wire_827,
fourFunc_wire_828,
fourFunc_wire_829,
fourFunc_wire_830,
fourFunc_wire_831,
fourFunc_wire_832,
fourFunc_wire_833,
fourFunc_wire_834,
fourFunc_wire_835,
fourFunc_wire_836,
fourFunc_wire_837,
fourFunc_wire_838,
fourFunc_wire_839,
fourFunc_wire_840,
fourFunc_wire_841,
fourFunc_wire_842,
fourFunc_wire_843,
fourFunc_wire_844,
fourFunc_wire_845,
fourFunc_wire_846,
fourFunc_wire_847,
fourFunc_wire_848,
fourFunc_wire_849,
fourFunc_wire_850,
fourFunc_wire_851,
fourFunc_wire_852,
fourFunc_wire_853,
fourFunc_wire_854,
fourFunc_wire_855,
fourFunc_wire_856,
fourFunc_wire_857,
fourFunc_wire_858,
fourFunc_wire_859,
fourFunc_wire_860,
fourFunc_wire_861,
fourFunc_wire_862,
fourFunc_wire_863,
fourFunc_wire_864,
fourFunc_wire_865,
fourFunc_wire_866,
fourFunc_wire_867,
fourFunc_wire_868,
fourFunc_wire_869,
fourFunc_wire_870,
fourFunc_wire_871,
fourFunc_wire_54_0,
fourFunc_wire_54_1,
fourFunc_wire_54_2,
fourFunc_wire_57_0,
fourFunc_wire_57_1,
fourFunc_wire_57_2,
fourFunc_wire_62_0,
fourFunc_wire_62_1,
fourFunc_wire_62_2,
fourFunc_wire_67_0,
fourFunc_wire_67_1,
fourFunc_wire_67_2,
fourFunc_wire_72_0,
fourFunc_wire_72_1,
fourFunc_wire_72_2,
fourFunc_wire_77_0,
fourFunc_wire_77_1,
fourFunc_wire_77_2,
fourFunc_wire_87_0,
fourFunc_wire_87_1,
fourFunc_wire_87_2,
fourFunc_wire_92_0,
fourFunc_wire_92_1,
fourFunc_wire_92_2,
fourFunc_wire_96_0,
fourFunc_wire_96_1,
fourFunc_wire_96_2,
fourFunc_wire_100_0,
fourFunc_wire_100_1,
fourFunc_wire_100_2,
fourFunc_wire_104_0,
fourFunc_wire_104_1,
fourFunc_wire_104_2,
fourFunc_wire_108_0,
fourFunc_wire_108_1,
fourFunc_wire_108_2,
fourFunc_wire_116_0,
fourFunc_wire_116_1,
fourFunc_wire_116_2,
fourFunc_wire_121_0,
fourFunc_wire_121_1,
fourFunc_wire_121_2,
fourFunc_wire_125_0,
fourFunc_wire_125_1,
fourFunc_wire_125_2,
fourFunc_wire_129_0,
fourFunc_wire_129_1,
fourFunc_wire_129_2,
fourFunc_wire_133_0,
fourFunc_wire_133_1,
fourFunc_wire_133_2,
fourFunc_wire_137_0,
fourFunc_wire_137_1,
fourFunc_wire_137_2,
fourFunc_wire_145_0,
fourFunc_wire_145_1,
fourFunc_wire_145_2,
fourFunc_wire_150_0,
fourFunc_wire_150_1,
fourFunc_wire_150_2,
fourFunc_wire_154_0,
fourFunc_wire_154_1,
fourFunc_wire_154_2,
fourFunc_wire_158_0,
fourFunc_wire_158_1,
fourFunc_wire_158_2,
fourFunc_wire_162_0,
fourFunc_wire_162_1,
fourFunc_wire_162_2,
fourFunc_wire_166_0,
fourFunc_wire_166_1,
fourFunc_wire_166_2,
fourFunc_wire_174_0,
fourFunc_wire_174_1,
fourFunc_wire_174_2,
fourFunc_wire_179_0,
fourFunc_wire_179_1,
fourFunc_wire_179_2,
fourFunc_wire_183_0,
fourFunc_wire_183_1,
fourFunc_wire_183_2,
fourFunc_wire_187_0,
fourFunc_wire_187_1,
fourFunc_wire_187_2,
fourFunc_wire_191_0,
fourFunc_wire_191_1,
fourFunc_wire_191_2,
fourFunc_wire_195_0,
fourFunc_wire_195_1,
fourFunc_wire_195_2,
fourFunc_wire_203_0,
fourFunc_wire_203_1,
fourFunc_wire_203_2,
fourFunc_wire_208_0,
fourFunc_wire_208_1,
fourFunc_wire_208_2,
fourFunc_wire_212_0,
fourFunc_wire_212_1,
fourFunc_wire_212_2,
fourFunc_wire_216_0,
fourFunc_wire_216_1,
fourFunc_wire_216_2,
fourFunc_wire_220_0,
fourFunc_wire_220_1,
fourFunc_wire_220_2,
fourFunc_wire_224_0,
fourFunc_wire_224_1,
fourFunc_wire_224_2,
fourFunc_wire_84_0,
fourFunc_wire_84_1,
fourFunc_wire_79_0,
fourFunc_wire_79_1,
fourFunc_wire_74_0,
fourFunc_wire_74_1,
fourFunc_wire_69_0,
fourFunc_wire_69_1,
fourFunc_wire_64_0,
fourFunc_wire_64_1,
fourFunc_wire_59_0,
fourFunc_wire_59_1,
fourFunc_wire_56_0,
fourFunc_wire_56_1,
fourFunc_wire_91_0,
fourFunc_wire_91_1,
fourFunc_wire_91_2,
fourFunc_wire_114_0,
fourFunc_wire_114_1,
fourFunc_wire_110_0,
fourFunc_wire_110_1,
fourFunc_wire_106_0,
fourFunc_wire_106_1,
fourFunc_wire_102_0,
fourFunc_wire_102_1,
fourFunc_wire_98_0,
fourFunc_wire_98_1,
fourFunc_wire_94_0,
fourFunc_wire_94_1,
fourFunc_wire_89_0,
fourFunc_wire_89_1,
fourFunc_wire_120_0,
fourFunc_wire_120_1,
fourFunc_wire_120_2,
fourFunc_wire_143_0,
fourFunc_wire_143_1,
fourFunc_wire_139_0,
fourFunc_wire_139_1,
fourFunc_wire_135_0,
fourFunc_wire_135_1,
fourFunc_wire_131_0,
fourFunc_wire_131_1,
fourFunc_wire_127_0,
fourFunc_wire_127_1,
fourFunc_wire_123_0,
fourFunc_wire_123_1,
fourFunc_wire_118_0,
fourFunc_wire_118_1,
fourFunc_wire_149_0,
fourFunc_wire_149_1,
fourFunc_wire_149_2,
fourFunc_wire_172_0,
fourFunc_wire_172_1,
fourFunc_wire_168_0,
fourFunc_wire_168_1,
fourFunc_wire_164_0,
fourFunc_wire_164_1,
fourFunc_wire_160_0,
fourFunc_wire_160_1,
fourFunc_wire_156_0,
fourFunc_wire_156_1,
fourFunc_wire_152_0,
fourFunc_wire_152_1,
fourFunc_wire_147_0,
fourFunc_wire_147_1,
fourFunc_wire_178_0,
fourFunc_wire_178_1,
fourFunc_wire_178_2,
fourFunc_wire_201_0,
fourFunc_wire_201_1,
fourFunc_wire_197_0,
fourFunc_wire_197_1,
fourFunc_wire_193_0,
fourFunc_wire_193_1,
fourFunc_wire_189_0,
fourFunc_wire_189_1,
fourFunc_wire_185_0,
fourFunc_wire_185_1,
fourFunc_wire_181_0,
fourFunc_wire_181_1,
fourFunc_wire_176_0,
fourFunc_wire_176_1,
fourFunc_wire_207_0,
fourFunc_wire_207_1,
fourFunc_wire_207_2,
fourFunc_wire_230_0,
fourFunc_wire_230_1,
fourFunc_wire_226_0,
fourFunc_wire_226_1,
fourFunc_wire_222_0,
fourFunc_wire_222_1,
fourFunc_wire_218_0,
fourFunc_wire_218_1,
fourFunc_wire_214_0,
fourFunc_wire_214_1,
fourFunc_wire_210_0,
fourFunc_wire_210_1,
fourFunc_wire_205_0,
fourFunc_wire_205_1,
fourFunc_wire_236_0,
fourFunc_wire_236_1,
fourFunc_wire_236_2,
fourFunc_wire_259_0,
fourFunc_wire_259_1,
fourFunc_wire_255_0,
fourFunc_wire_255_1,
fourFunc_wire_251_0,
fourFunc_wire_251_1,
fourFunc_wire_247_0,
fourFunc_wire_247_1,
fourFunc_wire_243_0,
fourFunc_wire_243_1,
fourFunc_wire_239_0,
fourFunc_wire_239_1,
fourFunc_wire_234_0,
fourFunc_wire_234_1,
fourFunc_wire_61_0,
fourFunc_wire_61_1,
fourFunc_wire_61_2,
fourFunc_wire_66_0,
fourFunc_wire_66_1,
fourFunc_wire_66_2,
fourFunc_wire_71_0,
fourFunc_wire_71_1,
fourFunc_wire_71_2,
fourFunc_wire_76_0,
fourFunc_wire_76_1,
fourFunc_wire_76_2,
fourFunc_wire_81_0,
fourFunc_wire_81_1,
fourFunc_wire_81_2,
fourFunc_wire_86_0,
fourFunc_wire_86_1,
fourFunc_wire_86_2,
fourFunc_wire_261_0,
fourFunc_wire_261_1,
fourFunc_wire_60_0,
fourFunc_wire_60_1,
fourFunc_wire_60_2,
fourFunc_wire_65_0,
fourFunc_wire_65_1,
fourFunc_wire_65_2,
fourFunc_wire_70_0,
fourFunc_wire_70_1,
fourFunc_wire_70_2,
fourFunc_wire_75_0,
fourFunc_wire_75_1,
fourFunc_wire_75_2,
fourFunc_wire_80_0,
fourFunc_wire_80_1,
fourFunc_wire_80_2,
fourFunc_wire_85_0,
fourFunc_wire_85_1,
fourFunc_wire_85_2,
fourFunc_wire_90_0,
fourFunc_wire_90_1,
fourFunc_wire_90_2,
fourFunc_wire_95_0,
fourFunc_wire_95_1,
fourFunc_wire_95_2,
fourFunc_wire_99_0,
fourFunc_wire_99_1,
fourFunc_wire_99_2,
fourFunc_wire_103_0,
fourFunc_wire_103_1,
fourFunc_wire_103_2,
fourFunc_wire_107_0,
fourFunc_wire_107_1,
fourFunc_wire_107_2,
fourFunc_wire_111_0,
fourFunc_wire_111_1,
fourFunc_wire_111_2,
fourFunc_wire_115_0,
fourFunc_wire_115_1,
fourFunc_wire_115_2,
fourFunc_wire_119_0,
fourFunc_wire_119_1,
fourFunc_wire_119_2,
fourFunc_wire_124_0,
fourFunc_wire_124_1,
fourFunc_wire_124_2,
fourFunc_wire_128_0,
fourFunc_wire_128_1,
fourFunc_wire_128_2,
fourFunc_wire_132_0,
fourFunc_wire_132_1,
fourFunc_wire_132_2,
fourFunc_wire_136_0,
fourFunc_wire_136_1,
fourFunc_wire_136_2,
fourFunc_wire_140_0,
fourFunc_wire_140_1,
fourFunc_wire_140_2,
fourFunc_wire_144_0,
fourFunc_wire_144_1,
fourFunc_wire_144_2,
fourFunc_wire_148_0,
fourFunc_wire_148_1,
fourFunc_wire_148_2,
fourFunc_wire_153_0,
fourFunc_wire_153_1,
fourFunc_wire_153_2,
fourFunc_wire_157_0,
fourFunc_wire_157_1,
fourFunc_wire_157_2,
fourFunc_wire_161_0,
fourFunc_wire_161_1,
fourFunc_wire_161_2,
fourFunc_wire_165_0,
fourFunc_wire_165_1,
fourFunc_wire_165_2,
fourFunc_wire_169_0,
fourFunc_wire_169_1,
fourFunc_wire_169_2,
fourFunc_wire_173_0,
fourFunc_wire_173_1,
fourFunc_wire_173_2,
fourFunc_wire_177_0,
fourFunc_wire_177_1,
fourFunc_wire_177_2,
fourFunc_wire_182_0,
fourFunc_wire_182_1,
fourFunc_wire_182_2,
fourFunc_wire_186_0,
fourFunc_wire_186_1,
fourFunc_wire_186_2,
fourFunc_wire_190_0,
fourFunc_wire_190_1,
fourFunc_wire_190_2,
fourFunc_wire_194_0,
fourFunc_wire_194_1,
fourFunc_wire_194_2,
fourFunc_wire_198_0,
fourFunc_wire_198_1,
fourFunc_wire_198_2,
fourFunc_wire_202_0,
fourFunc_wire_202_1,
fourFunc_wire_202_2,
fourFunc_wire_206_0,
fourFunc_wire_206_1,
fourFunc_wire_206_2,
fourFunc_wire_211_0,
fourFunc_wire_211_1,
fourFunc_wire_211_2,
fourFunc_wire_215_0,
fourFunc_wire_215_1,
fourFunc_wire_215_2,
fourFunc_wire_219_0,
fourFunc_wire_219_1,
fourFunc_wire_219_2,
fourFunc_wire_223_0,
fourFunc_wire_223_1,
fourFunc_wire_223_2,
fourFunc_wire_227_0,
fourFunc_wire_227_1,
fourFunc_wire_227_2,
fourFunc_wire_231_0,
fourFunc_wire_231_1,
fourFunc_wire_231_2,
fourFunc_wire_235_0,
fourFunc_wire_235_1,
fourFunc_wire_235_2,
fourFunc_wire_240_0,
fourFunc_wire_240_1,
fourFunc_wire_240_2,
fourFunc_wire_244_0,
fourFunc_wire_244_1,
fourFunc_wire_244_2,
fourFunc_wire_248_0,
fourFunc_wire_248_1,
fourFunc_wire_248_2,
fourFunc_wire_252_0,
fourFunc_wire_252_1,
fourFunc_wire_252_2,
fourFunc_wire_256_0,
fourFunc_wire_256_1,
fourFunc_wire_256_2,
fourFunc_wire_260_0,
fourFunc_wire_260_1,
fourFunc_wire_260_2,
fourFunc_wire_502_0,
fourFunc_wire_502_1,
fourFunc_wire_499_0,
fourFunc_wire_499_1,
fourFunc_wire_496_0,
fourFunc_wire_496_1,
fourFunc_wire_493_0,
fourFunc_wire_493_1,
fourFunc_wire_490_0,
fourFunc_wire_490_1,
fourFunc_wire_487_0,
fourFunc_wire_487_1,
fourFunc_wire_484_0,
fourFunc_wire_484_1,
fourFunc_wire_479_0,
fourFunc_wire_479_1,
fourFunc_wire_475_0,
fourFunc_wire_475_1,
fourFunc_wire_471_0,
fourFunc_wire_471_1,
fourFunc_wire_467_0,
fourFunc_wire_467_1,
fourFunc_wire_463_0,
fourFunc_wire_463_1,
fourFunc_wire_459_0,
fourFunc_wire_459_1,
fourFunc_wire_455_0,
fourFunc_wire_455_1,
fourFunc_wire_451_0,
fourFunc_wire_451_1,
fourFunc_wire_448_0,
fourFunc_wire_448_1,
fourFunc_wire_448_2,
fourFunc_wire_563_0,
fourFunc_wire_563_1,
fourFunc_wire_563_2,
fourFunc_wire_563_3,
fourFunc_wire_563_4,
fourFunc_wire_563_5,
fourFunc_wire_563_6,
fourFunc_wire_563_7,
fourFunc_wire_563_8,
fourFunc_wire_563_9,
fourFunc_wire_563_10,
fourFunc_wire_563_11,
fourFunc_wire_563_12,
fourFunc_wire_563_13,
fourFunc_wire_563_14,
fourFunc_wire_563_15,
fourFunc_wire_563_16,
fourFunc_wire_563_17,
fourFunc_wire_563_18,
fourFunc_wire_563_19,
fourFunc_wire_563_20,
fourFunc_wire_563_21,
fourFunc_wire_11_0,
fourFunc_wire_11_1,
fourFunc_wire_11_2,
fourFunc_wire_11_3,
fourFunc_wire_11_4,
fourFunc_wire_11_5,
fourFunc_wire_11_6,
fourFunc_wire_11_7,
fourFunc_wire_11_8,
fourFunc_wire_11_9,
fourFunc_wire_11_10,
fourFunc_wire_11_11,
fourFunc_wire_11_12,
fourFunc_wire_11_13,
fourFunc_wire_3_0,
fourFunc_wire_3_1,
fourFunc_wire_3_2,
fourFunc_wire_3_3,
fourFunc_wire_3_4,
fourFunc_wire_3_5,
fourFunc_wire_3_6,
fourFunc_wire_3_7,
fourFunc_wire_3_8,
fourFunc_wire_3_9,
fourFunc_wire_3_10,
fourFunc_wire_3_11,
fourFunc_wire_3_12,
fourFunc_wire_3_13,
fourFunc_wire_2_0,
fourFunc_wire_2_1,
fourFunc_wire_2_2,
fourFunc_wire_2_3,
fourFunc_wire_2_4,
fourFunc_wire_2_5,
fourFunc_wire_2_6,
fourFunc_wire_2_7,
fourFunc_wire_2_8,
fourFunc_wire_2_9,
fourFunc_wire_2_10,
fourFunc_wire_2_11,
fourFunc_wire_2_12,
fourFunc_wire_2_13,
fourFunc_wire_2_14,
fourFunc_wire_2_15,
fourFunc_wire_2_16,
fourFunc_wire_2_17,
fourFunc_wire_2_18,
fourFunc_wire_564_0,
fourFunc_wire_564_1,
fourFunc_wire_565_0,
fourFunc_wire_565_1,
fourFunc_wire_566_0,
fourFunc_wire_566_1,
fourFunc_wire_567_0,
fourFunc_wire_567_1,
fourFunc_wire_568_0,
fourFunc_wire_568_1,
fourFunc_wire_569_0,
fourFunc_wire_569_1,
fourFunc_wire_570_0,
fourFunc_wire_570_1,
fourFunc_wire_571_0,
fourFunc_wire_571_1,
fourFunc_wire_422_0,
fourFunc_wire_422_1,
fourFunc_wire_422_2,
fourFunc_wire_422_3,
fourFunc_wire_422_4,
fourFunc_wire_422_5,
fourFunc_wire_422_6,
fourFunc_wire_422_7,
fourFunc_wire_422_8,
fourFunc_wire_422_9,
fourFunc_wire_422_10,
fourFunc_wire_422_11,
fourFunc_wire_430_0,
fourFunc_wire_430_1,
fourFunc_wire_430_2,
fourFunc_wire_430_3,
fourFunc_wire_430_4,
fourFunc_wire_430_5,
fourFunc_wire_430_6,
fourFunc_wire_430_7,
fourFunc_wire_430_8,
fourFunc_wire_430_9,
fourFunc_wire_430_10,
fourFunc_wire_430_11,
fourFunc_wire_430_12,
fourFunc_wire_430_13,
fourFunc_wire_430_14,
fourFunc_wire_432_0,
fourFunc_wire_432_1,
fourFunc_wire_432_2,
fourFunc_wire_432_3,
fourFunc_wire_432_4,
fourFunc_wire_432_5,
fourFunc_wire_432_6,
fourFunc_wire_432_7,
fourFunc_wire_432_8,
fourFunc_wire_432_9,
fourFunc_wire_432_10,
fourFunc_wire_432_11,
fourFunc_wire_432_12,
fourFunc_wire_432_13,
fourFunc_wire_432_14,
fourFunc_wire_433_0,
fourFunc_wire_433_1,
fourFunc_wire_433_2,
fourFunc_wire_433_3,
fourFunc_wire_433_4,
fourFunc_wire_433_5,
fourFunc_wire_433_6,
fourFunc_wire_433_7,
fourFunc_wire_433_8,
fourFunc_wire_433_9,
fourFunc_wire_433_10,
fourFunc_wire_433_11,
fourFunc_wire_433_12,
fourFunc_wire_433_13,
fourFunc_wire_433_14,
fourFunc_wire_434_0,
fourFunc_wire_434_1,
fourFunc_wire_434_2,
fourFunc_wire_434_3,
fourFunc_wire_434_4,
fourFunc_wire_434_5,
fourFunc_wire_434_6,
fourFunc_wire_434_7,
fourFunc_wire_434_8,
fourFunc_wire_434_9,
fourFunc_wire_434_10,
fourFunc_wire_434_11,
fourFunc_wire_434_12,
fourFunc_wire_434_13,
fourFunc_wire_434_14,
fourFunc_wire_435_0,
fourFunc_wire_435_1,
fourFunc_wire_435_2,
fourFunc_wire_435_3,
fourFunc_wire_435_4,
fourFunc_wire_435_5,
fourFunc_wire_435_6,
fourFunc_wire_435_7,
fourFunc_wire_435_8,
fourFunc_wire_435_9,
fourFunc_wire_435_10,
fourFunc_wire_435_11,
fourFunc_wire_435_12,
fourFunc_wire_435_13,
fourFunc_wire_435_14,
fourFunc_wire_436_0,
fourFunc_wire_436_1,
fourFunc_wire_436_2,
fourFunc_wire_436_3,
fourFunc_wire_436_4,
fourFunc_wire_436_5,
fourFunc_wire_436_6,
fourFunc_wire_436_7,
fourFunc_wire_436_8,
fourFunc_wire_436_9,
fourFunc_wire_436_10,
fourFunc_wire_436_11,
fourFunc_wire_436_12,
fourFunc_wire_436_13,
fourFunc_wire_436_14,
fourFunc_wire_437_0,
fourFunc_wire_437_1,
fourFunc_wire_437_2,
fourFunc_wire_437_3,
fourFunc_wire_437_4,
fourFunc_wire_437_5,
fourFunc_wire_437_6,
fourFunc_wire_437_7,
fourFunc_wire_437_8,
fourFunc_wire_437_9,
fourFunc_wire_437_10,
fourFunc_wire_437_11,
fourFunc_wire_437_12,
fourFunc_wire_437_13,
fourFunc_wire_437_14,
fourFunc_wire_442_0,
fourFunc_wire_442_1,
fourFunc_wire_442_2,
fourFunc_wire_442_3,
fourFunc_wire_442_4,
fourFunc_wire_442_5,
fourFunc_wire_476_0,
fourFunc_wire_476_1,
fourFunc_wire_476_2,
fourFunc_wire_476_3,
fourFunc_wire_476_4,
fourFunc_wire_476_5,
fourFunc_wire_476_6,
fourFunc_wire_476_7,
fourFunc_wire_472_0,
fourFunc_wire_472_1,
fourFunc_wire_472_2,
fourFunc_wire_472_3,
fourFunc_wire_472_4,
fourFunc_wire_472_5,
fourFunc_wire_472_6,
fourFunc_wire_472_7,
fourFunc_wire_468_0,
fourFunc_wire_468_1,
fourFunc_wire_468_2,
fourFunc_wire_468_3,
fourFunc_wire_468_4,
fourFunc_wire_468_5,
fourFunc_wire_468_6,
fourFunc_wire_468_7,
fourFunc_wire_464_0,
fourFunc_wire_464_1,
fourFunc_wire_464_2,
fourFunc_wire_464_3,
fourFunc_wire_464_4,
fourFunc_wire_464_5,
fourFunc_wire_464_6,
fourFunc_wire_464_7,
fourFunc_wire_460_0,
fourFunc_wire_460_1,
fourFunc_wire_460_2,
fourFunc_wire_460_3,
fourFunc_wire_460_4,
fourFunc_wire_460_5,
fourFunc_wire_460_6,
fourFunc_wire_460_7,
fourFunc_wire_456_0,
fourFunc_wire_456_1,
fourFunc_wire_456_2,
fourFunc_wire_456_3,
fourFunc_wire_456_4,
fourFunc_wire_456_5,
fourFunc_wire_456_6,
fourFunc_wire_456_7,
fourFunc_wire_452_0,
fourFunc_wire_452_1,
fourFunc_wire_452_2,
fourFunc_wire_452_3,
fourFunc_wire_452_4,
fourFunc_wire_452_5,
fourFunc_wire_452_6,
fourFunc_wire_452_7,
fourFunc_wire_447_0,
fourFunc_wire_447_1,
fourFunc_wire_447_2,
fourFunc_wire_447_3,
fourFunc_wire_447_4,
fourFunc_wire_447_5,
fourFunc_wire_447_6,
fourFunc_wire_444_0,
fourFunc_wire_444_1,
fourFunc_wire_444_2,
fourFunc_wire_444_3,
fourFunc_wire_594_0,
fourFunc_wire_594_1,
fourFunc_wire_600_0,
fourFunc_wire_600_1,
fourFunc_wire_600_2,
fourFunc_wire_600_3,
fourFunc_wire_601_0,
fourFunc_wire_601_1,
fourFunc_wire_601_2,
fourFunc_wire_601_3,
fourFunc_wire_601_4,
fourFunc_wire_602_0,
fourFunc_wire_602_1,
fourFunc_wire_602_2,
fourFunc_wire_598_0,
fourFunc_wire_598_1,
fourFunc_wire_598_2,
fourFunc_wire_598_3,
fourFunc_wire_598_4,
fourFunc_wire_598_5,
fourFunc_wire_598_6,
fourFunc_wire_598_7,
fourFunc_wire_598_8,
fourFunc_wire_598_9,
fourFunc_wire_598_10,
fourFunc_wire_598_11,
fourFunc_wire_598_12,
fourFunc_wire_598_13,
fourFunc_wire_598_14,
fourFunc_wire_598_15,
fourFunc_wire_598_16,
fourFunc_wire_598_17,
fourFunc_wire_598_18,
fourFunc_wire_598_19,
fourFunc_wire_593_0,
fourFunc_wire_593_1,
fourFunc_wire_593_2,
fourFunc_wire_593_3,
fourFunc_wire_593_4,
fourFunc_wire_611_0,
fourFunc_wire_611_1,
fourFunc_wire_611_2,
fourFunc_wire_611_3,
fourFunc_wire_611_4,
fourFunc_wire_611_5,
fourFunc_wire_611_6,
fourFunc_wire_611_7,
fourFunc_wire_611_8,
fourFunc_wire_611_9,
fourFunc_wire_611_10,
fourFunc_wire_611_11,
fourFunc_wire_611_12,
fourFunc_wire_611_13,
fourFunc_wire_611_14,
fourFunc_wire_611_15,
fourFunc_wire_611_16,
fourFunc_wire_611_17,
fourFunc_wire_611_18,
fourFunc_wire_611_19,
fourFunc_wire_611_20,
fourFunc_wire_611_21,
fourFunc_wire_611_22,
fourFunc_wire_611_23,
fourFunc_wire_611_24,
fourFunc_wire_611_25,
fourFunc_wire_611_26,
fourFunc_wire_611_27,
fourFunc_wire_611_28,
fourFunc_wire_611_29,
fourFunc_wire_611_30,
fourFunc_wire_611_31,
fourFunc_wire_612_0,
fourFunc_wire_612_1,
fourFunc_wire_618_0,
fourFunc_wire_618_1,
fourFunc_wire_622_0,
fourFunc_wire_622_1,
fourFunc_wire_622_2,
fourFunc_wire_621_0,
fourFunc_wire_621_1,
fourFunc_wire_621_2,
fourFunc_wire_621_3,
fourFunc_wire_621_4,
fourFunc_wire_621_5,
fourFunc_wire_621_6,
fourFunc_wire_621_7,
fourFunc_wire_621_8,
fourFunc_wire_621_9,
fourFunc_wire_621_10,
fourFunc_wire_621_11,
fourFunc_wire_617_0,
fourFunc_wire_617_1,
fourFunc_wire_617_2,
fourFunc_wire_617_3,
fourFunc_wire_617_4,
fourFunc_wire_617_5,
fourFunc_wire_617_6,
fourFunc_wire_617_7,
fourFunc_wire_617_8,
fourFunc_wire_617_9,
fourFunc_wire_617_10,
fourFunc_wire_617_11,
fourFunc_wire_617_12,
fourFunc_wire_617_13,
fourFunc_wire_617_14,
fourFunc_wire_617_15,
fourFunc_wire_617_16,
fourFunc_wire_617_17,
fourFunc_wire_617_18,
fourFunc_wire_617_19,
fourFunc_wire_617_20,
fourFunc_wire_617_21,
fourFunc_wire_617_22,
fourFunc_wire_617_23,
fourFunc_wire_617_24,
fourFunc_wire_617_25,
fourFunc_wire_617_26,
fourFunc_wire_617_27,
fourFunc_wire_617_28,
fourFunc_wire_617_29,
fourFunc_wire_617_30,
fourFunc_wire_617_31,
fourFunc_wire_617_32,
fourFunc_wire_617_33,
fourFunc_wire_617_34,
fourFunc_wire_617_35,
fourFunc_wire_617_36,
fourFunc_wire_617_37,
fourFunc_wire_617_38,
fourFunc_wire_617_39,
fourFunc_wire_659_0,
fourFunc_wire_659_1,
fourFunc_wire_659_2,
fourFunc_wire_659_3,
fourFunc_wire_659_4,
fourFunc_wire_659_5,
fourFunc_wire_659_6,
fourFunc_wire_659_7,
fourFunc_wire_659_8,
fourFunc_wire_659_9,
fourFunc_wire_659_10,
fourFunc_wire_431_0,
fourFunc_wire_431_1,
fourFunc_wire_431_2,
fourFunc_wire_431_3,
fourFunc_wire_431_4,
fourFunc_wire_431_5,
fourFunc_wire_431_6,
fourFunc_wire_429_0,
fourFunc_wire_429_1,
fourFunc_wire_429_2,
fourFunc_wire_429_3,
fourFunc_wire_429_4,
fourFunc_wire_429_5,
fourFunc_wire_429_6,
fourFunc_wire_429_7,
fourFunc_wire_428_0,
fourFunc_wire_428_1,
fourFunc_wire_428_2,
fourFunc_wire_428_3,
fourFunc_wire_428_4,
fourFunc_wire_428_5,
fourFunc_wire_428_6,
fourFunc_wire_428_7,
fourFunc_wire_427_0,
fourFunc_wire_427_1,
fourFunc_wire_427_2,
fourFunc_wire_427_3,
fourFunc_wire_427_4,
fourFunc_wire_427_5,
fourFunc_wire_427_6,
fourFunc_wire_427_7,
fourFunc_wire_426_0,
fourFunc_wire_426_1,
fourFunc_wire_426_2,
fourFunc_wire_426_3,
fourFunc_wire_426_4,
fourFunc_wire_426_5,
fourFunc_wire_426_6,
fourFunc_wire_426_7,
fourFunc_wire_425_0,
fourFunc_wire_425_1,
fourFunc_wire_425_2,
fourFunc_wire_425_3,
fourFunc_wire_425_4,
fourFunc_wire_425_5,
fourFunc_wire_425_6,
fourFunc_wire_425_7,
fourFunc_wire_424_0,
fourFunc_wire_424_1,
fourFunc_wire_424_2,
fourFunc_wire_424_3,
fourFunc_wire_424_4,
fourFunc_wire_424_5,
fourFunc_wire_424_6,
fourFunc_wire_424_7,
fourFunc_wire_423_0,
fourFunc_wire_423_1,
fourFunc_wire_423_2,
fourFunc_wire_423_3,
fourFunc_wire_423_4,
fourFunc_wire_423_5,
fourFunc_wire_423_6,
fourFunc_wire_423_7,
fourFunc_wire_733_0,
fourFunc_wire_733_1,
fourFunc_wire_733_2,
fourFunc_wire_733_3,
fourFunc_wire_733_4,
fourFunc_wire_733_5,
fourFunc_wire_733_6,
fourFunc_wire_733_7,
fourFunc_wire_733_8,
fourFunc_wire_7_0,
fourFunc_wire_7_1,
fourFunc_wire_7_2,
fourFunc_wire_7_3,
fourFunc_wire_7_4,
fourFunc_wire_7_5,
fourFunc_wire_7_6,
fourFunc_wire_7_7,
fourFunc_wire_7_8,
fourFunc_wire_7_9,
fourFunc_wire_7_10,
fourFunc_wire_7_11,
fourFunc_wire_7_12,
fourFunc_wire_7_13,
fourFunc_wire_7_14,
fourFunc_wire_7_15,
fourFunc_wire_7_16,
fourFunc_wire_7_17,
fourFunc_wire_7_18,
fourFunc_wire_7_19,
fourFunc_wire_7_20,
fourFunc_wire_7_21,
fourFunc_wire_7_22,
fourFunc_wire_7_23,
fourFunc_wire_7_24,
fourFunc_wire_7_25,
fourFunc_wire_7_26,
fourFunc_wire_7_27,
fourFunc_wire_7_28,
fourFunc_wire_7_29,
fourFunc_wire_7_30,
fourFunc_wire_7_31,
fourFunc_wire_610_0,
fourFunc_wire_610_1,
fourFunc_wire_610_2,
fourFunc_wire_610_3,
fourFunc_wire_610_4,
fourFunc_wire_610_5,
fourFunc_wire_650_0,
fourFunc_wire_650_1,
fourFunc_wire_650_2,
fourFunc_wire_637_0,
fourFunc_wire_637_1,
fourFunc_wire_637_2,
fourFunc_wire_639_0,
fourFunc_wire_639_1,
fourFunc_wire_639_2,
fourFunc_wire_641_0,
fourFunc_wire_641_1,
fourFunc_wire_641_2,
fourFunc_wire_635_0,
fourFunc_wire_635_1,
fourFunc_wire_635_2,
fourFunc_wire_643_0,
fourFunc_wire_643_1,
fourFunc_wire_643_2,
fourFunc_wire_645_0,
fourFunc_wire_645_1,
fourFunc_wire_645_2,
fourFunc_wire_647_0,
fourFunc_wire_647_1,
fourFunc_wire_647_2,
fourFunc_wire_649_0,
fourFunc_wire_649_1,
fourFunc_wire_649_2,
NOT_intermediateXXXwire_735_0,
NOT_intermediateXXXwire_735_1,
NOT_intermediateXXXwire_739_0,
NOT_intermediateXXXwire_739_1,
NOT_intermediateXXXwire_739_2,
NOT_intermediateXXXwire_739_3,
NOT_intermediateXXXwire_739_4,
NOT_intermediateXXXwire_739_5,
NOT_intermediateXXXwire_739_6,
NOT_intermediateXXXwire_739_7,
NOT_intermediateXXXwire_963_0,
NOT_intermediateXXXwire_963_1,
NOT_intermediateXXXwire_963_2,
NOT_intermediateXXXwire_963_3,
NOT_intermediateXXXwire_963_4,
NOT_intermediateXXXwire_963_5,
NOT_intermediateXXXwire_963_6,
NOT_intermediateXXXwire_963_7,
NOT_intermediateXXXwire_834_0,
NOT_intermediateXXXwire_834_1,
NOT_intermediateXXXwire_834_2,
NOT_intermediateXXXwire_834_3,
NOT_intermediateXXXwire_834_4,
NOT_intermediateXXXwire_834_5,
NOT_intermediateXXXwire_834_6,
NOT_intermediateXXXwire_834_7,
NOT_intermediateXXXwire_834_8,
NOT_intermediateXXXwire_834_9,
clk_net_0,
rst_net_0,
start_net_0,
busy_net_0 ;
//PPI
/* fourFunc_wire_563,
fourFunc_wire_11,
fourFunc_wire_3,
fourFunc_wire_2,
fourFunc_wire_564,
fourFunc_wire_565,
fourFunc_wire_566,
fourFunc_wire_567,
fourFunc_wire_568,
fourFunc_wire_569,
fourFunc_wire_570,
fourFunc_wire_571,
fourFunc_wire_422,
fourFunc_wire_430,
fourFunc_wire_432,
fourFunc_wire_433,
fourFunc_wire_434,
fourFunc_wire_435,
fourFunc_wire_436,
fourFunc_wire_437,
fourFunc_wire_442,
fourFunc_wire_476,
fourFunc_wire_472,
fourFunc_wire_468,
fourFunc_wire_464,
fourFunc_wire_460,
fourFunc_wire_456,
fourFunc_wire_452,
fourFunc_wire_447,
fourFunc_wire_444,
fourFunc_wire_604,
fourFunc_wire_600,
fourFunc_wire_601,
fourFunc_wire_602,
fourFunc_wire_598,
fourFunc_wire_593,
fourFunc_wire_611,
NOT_intermediateXXXwire_721_AND_intermediateXXXwire_718_OR_intermediateXXXwire_721_AND_intermediateXXXwire_719,
NOT_intermediateXXXwire_731_AND_intermediateXXXwire_61_OR_intermediateXXXwire_731_AND_intermediateXXXwire_727,
NOT_intermediateXXXwire_735_AND_intermediateXXXwire_63_OR_intermediateXXXwire_735_AND_intermediateXXXwire_737,
NOT_intermediateXXXwire_735_AND_intermediateXXXwire_62_OR_intermediateXXXwire_735_AND_intermediateXXXwire_733,
NOT_intermediateXXXwire_739_AND_intermediateXXXwire_796_OR_intermediateXXXwire_739_AND_intermediateXXXwire_797,
NOT_intermediateXXXwire_739_AND_intermediateXXXwire_799_OR_intermediateXXXwire_739_AND_intermediateXXXwire_800,
NOT_intermediateXXXwire_739_AND_intermediateXXXwire_802_OR_intermediateXXXwire_739_AND_intermediateXXXwire_803,
NOT_intermediateXXXwire_739_AND_intermediateXXXwire_805_OR_intermediateXXXwire_739_AND_intermediateXXXwire_806,
NOT_intermediateXXXwire_739_AND_intermediateXXXwire_808_OR_intermediateXXXwire_739_AND_intermediateXXXwire_809,
NOT_intermediateXXXwire_739_AND_intermediateXXXwire_811_OR_intermediateXXXwire_739_AND_intermediateXXXwire_812,
NOT_intermediateXXXwire_739_AND_intermediateXXXwire_814_OR_intermediateXXXwire_739_AND_intermediateXXXwire_815,
NOT_intermediateXXXwire_739_AND_intermediateXXXwire_817_OR_intermediateXXXwire_739_AND_intermediateXXXwire_818,
NOT_intermediateXXXwire_963_AND_intermediateXXXwire_955_OR_intermediateXXXwire_963_AND_intermediateXXXwire_956,
NOT_intermediateXXXwire_963_AND_intermediateXXXwire_965_OR_intermediateXXXwire_963_AND_intermediateXXXwire_966,
NOT_intermediateXXXwire_963_AND_intermediateXXXwire_973_OR_intermediateXXXwire_963_AND_intermediateXXXwire_974,
NOT_intermediateXXXwire_963_AND_intermediateXXXwire_981_OR_intermediateXXXwire_963_AND_intermediateXXXwire_982,
NOT_intermediateXXXwire_963_AND_intermediateXXXwire_989_OR_intermediateXXXwire_963_AND_intermediateXXXwire_990,
NOT_intermediateXXXwire_963_AND_intermediateXXXwire_997_OR_intermediateXXXwire_963_AND_intermediateXXXwire_998,
NOT_intermediateXXXwire_963_AND_intermediateXXXwire_1005_OR_intermediateXXXwire_963_AND_intermediateXXXwire_1006,
NOT_intermediateXXXwire_963_AND_intermediateXXXwire_1013_OR_intermediateXXXwire_963_AND_intermediateXXXwire_1014,
NOT_intermediateXXXwire_834_AND_intermediateXXXwire_820_OR_intermediateXXXwire_834_AND_intermediateXXXwire_821,
NOT_intermediateXXXwire_834_AND_intermediateXXXwire_835_OR_intermediateXXXwire_834_AND_intermediateXXXwire_836,
NOT_intermediateXXXwire_834_AND_intermediateXXXwire_848_OR_intermediateXXXwire_834_AND_intermediateXXXwire_849,
NOT_intermediateXXXwire_834_AND_intermediateXXXwire_861_OR_intermediateXXXwire_834_AND_intermediateXXXwire_862,
NOT_intermediateXXXwire_834_AND_intermediateXXXwire_874_OR_intermediateXXXwire_834_AND_intermediateXXXwire_875,
NOT_intermediateXXXwire_834_AND_intermediateXXXwire_887_OR_intermediateXXXwire_834_AND_intermediateXXXwire_888,
NOT_intermediateXXXwire_834_AND_intermediateXXXwire_900_OR_intermediateXXXwire_834_AND_intermediateXXXwire_901,
NOT_intermediateXXXwire_834_AND_intermediateXXXwire_913_OR_intermediateXXXwire_834_AND_intermediateXXXwire_914,
NOT_intermediateXXXwire_834_AND_intermediateXXXwire_926_OR_intermediateXXXwire_834_AND_intermediateXXXwire_927,
NOT_intermediateXXXwire_834_AND_intermediateXXXwire_937_OR_intermediateXXXwire_834_AND_intermediateXXXwire_938,
fourFunc_wire_603,
fourFunc_wire_605,
fourFunc_wire_606,
fourFunc_wire_607,
fourFunc_wire_608,
fourFunc_wire_609,
fourFunc_wire_610	*/
/////////////////////////////////////
//PPO


//pin #(13) pin_0 ({clk, rst, start, func[0], func[1], x[0], x[1], x[2], x[3], x[4], x[5], x[6], x[7]}, {clk_net_0, rst_net_0, start_net_0, func_0, func_1, x_0, x_1, x_2, x_3, x_4, x_5, x_6, x_7});
pin #(50) pin_0 ({clk, rst, start, func[0], func[1], x[0], x[1], x[2], x[3], x[4], x[5], x[6], x[7],PPI0, PPI1, PPI2, PPI3, PPI4, PPI5, PPI6, PPI7, PPI8, PPI9, PPI10, PPI11, PPI12, PPI13, PPI14, PPI15, PPI16, PPI17, PPI18, PPI19, PPI20, PPI21, PPI22, PPI23, PPI24, PPI25, PPI26, PPI27, PPI28, PPI29, PPI30, PPI31, PPI32, PPI33, PPI34, PPI35, PPI36}, {clk_net_0, rst_net_0, start_net_0, func_0, func_1, x_0, x_1, x_2, x_3, x_4, x_5, x_6, x_7, fourFunc_wire_563, fourFunc_wire_11, fourFunc_wire_3, fourFunc_wire_2, fourFunc_wire_564, fourFunc_wire_565, fourFunc_wire_566, fourFunc_wire_567, fourFunc_wire_568, fourFunc_wire_569, fourFunc_wire_570, fourFunc_wire_571, fourFunc_wire_422, fourFunc_wire_430, fourFunc_wire_432, fourFunc_wire_433, fourFunc_wire_434, fourFunc_wire_435, fourFunc_wire_436, fourFunc_wire_437, fourFunc_wire_442, fourFunc_wire_476, fourFunc_wire_472, fourFunc_wire_468, fourFunc_wire_464, fourFunc_wire_460, fourFunc_wire_456, fourFunc_wire_452, fourFunc_wire_447, fourFunc_wire_444, fourFunc_wire_604, fourFunc_wire_600, fourFunc_wire_601, fourFunc_wire_602, fourFunc_wire_598, fourFunc_wire_593, fourFunc_wire_611});

/////////////////////////////////////
/////////////////////////////////////




//pout #(11) pout_0 ({busy_net_0, resultIPart_0, resultIPart_1, resultFPart_0, resultFPart_1, resultFPart_2, resultFPart_3, resultFPart_4, resultFPart_5, resultFPart_6, resultFPart_7}, {busy, resultIPart[0], resultIPart[1], resultFPart[0], resultFPart[1], resultFPart[2], resultFPart[3], resultFPart[4], resultFPart[5], resultFPart[6], resultFPart[7]});
pout #(48) pout_0 ({busy_net_0, resultIPart_0, resultIPart_1, resultFPart_0, resultFPart_1, resultFPart_2, resultFPart_3, resultFPart_4, resultFPart_5, resultFPart_6, resultFPart_7,  NOT_intermediateXXXwire_721_AND_intermediateXXXwire_718_OR_intermediateXXXwire_721_AND_intermediateXXXwire_719, NOT_intermediateXXXwire_731_AND_intermediateXXXwire_61_OR_intermediateXXXwire_731_AND_intermediateXXXwire_727, NOT_intermediateXXXwire_735_AND_intermediateXXXwire_63_OR_intermediateXXXwire_735_AND_intermediateXXXwire_737, NOT_intermediateXXXwire_735_AND_intermediateXXXwire_62_OR_intermediateXXXwire_735_AND_intermediateXXXwire_733, NOT_intermediateXXXwire_739_AND_intermediateXXXwire_796_OR_intermediateXXXwire_739_AND_intermediateXXXwire_797, NOT_intermediateXXXwire_739_AND_intermediateXXXwire_799_OR_intermediateXXXwire_739_AND_intermediateXXXwire_800, NOT_intermediateXXXwire_739_AND_intermediateXXXwire_802_OR_intermediateXXXwire_739_AND_intermediateXXXwire_803, NOT_intermediateXXXwire_739_AND_intermediateXXXwire_805_OR_intermediateXXXwire_739_AND_intermediateXXXwire_806, NOT_intermediateXXXwire_739_AND_intermediateXXXwire_808_OR_intermediateXXXwire_739_AND_intermediateXXXwire_809, NOT_intermediateXXXwire_739_AND_intermediateXXXwire_811_OR_intermediateXXXwire_739_AND_intermediateXXXwire_812, NOT_intermediateXXXwire_739_AND_intermediateXXXwire_814_OR_intermediateXXXwire_739_AND_intermediateXXXwire_815, NOT_intermediateXXXwire_739_AND_intermediateXXXwire_817_OR_intermediateXXXwire_739_AND_intermediateXXXwire_818, NOT_intermediateXXXwire_963_AND_intermediateXXXwire_955_OR_intermediateXXXwire_963_AND_intermediateXXXwire_956, NOT_intermediateXXXwire_963_AND_intermediateXXXwire_965_OR_intermediateXXXwire_963_AND_intermediateXXXwire_966, NOT_intermediateXXXwire_963_AND_intermediateXXXwire_973_OR_intermediateXXXwire_963_AND_intermediateXXXwire_974, NOT_intermediateXXXwire_963_AND_intermediateXXXwire_981_OR_intermediateXXXwire_963_AND_intermediateXXXwire_982, NOT_intermediateXXXwire_963_AND_intermediateXXXwire_989_OR_intermediateXXXwire_963_AND_intermediateXXXwire_990, NOT_intermediateXXXwire_963_AND_intermediateXXXwire_997_OR_intermediateXXXwire_963_AND_intermediateXXXwire_998, NOT_intermediateXXXwire_963_AND_intermediateXXXwire_1005_OR_intermediateXXXwire_963_AND_intermediateXXXwire_1006, NOT_intermediateXXXwire_963_AND_intermediateXXXwire_1013_OR_intermediateXXXwire_963_AND_intermediateXXXwire_1014, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_820_OR_intermediateXXXwire_834_AND_intermediateXXXwire_821, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_835_OR_intermediateXXXwire_834_AND_intermediateXXXwire_836, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_848_OR_intermediateXXXwire_834_AND_intermediateXXXwire_849, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_861_OR_intermediateXXXwire_834_AND_intermediateXXXwire_862, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_874_OR_intermediateXXXwire_834_AND_intermediateXXXwire_875, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_887_OR_intermediateXXXwire_834_AND_intermediateXXXwire_888, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_900_OR_intermediateXXXwire_834_AND_intermediateXXXwire_901, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_913_OR_intermediateXXXwire_834_AND_intermediateXXXwire_914, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_926_OR_intermediateXXXwire_834_AND_intermediateXXXwire_927, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_937_OR_intermediateXXXwire_834_AND_intermediateXXXwire_938, fourFunc_wire_603, fourFunc_wire_605, fourFunc_wire_606, fourFunc_wire_607, fourFunc_wire_608, fourFunc_wire_609, fourFunc_wire_610}, {busy, resultIPart[0], resultIPart[1], resultFPart[0], resultFPart[1], resultFPart[2], resultFPart[3], resultFPart[4], resultFPart[5], resultFPart[6], resultFPart[7], PPO0, PPO1, PPO2, PPO3, PPO4, PPO5, PPO6, PPO7, PPO8, PPO9, PPO10, PPO11, PPO12, PPO13, PPO14, PPO15, PPO16, PPO17, PPO18, PPO19, PPO20, PPO21, PPO22, PPO23, PPO24, PPO25, PPO26, PPO27, PPO28, PPO29, PPO30, PPO31, PPO32, PPO33, PPO34, PPO35, PPO36});




////////////////////////////
fanout_n #(3, 0, 0) FANOUT_1 (fourFunc_wire_54, {fourFunc_wire_54_0, fourFunc_wire_54_1, fourFunc_wire_54_2});
fanout_n #(3, 0, 0) FANOUT_2 (fourFunc_wire_57, {fourFunc_wire_57_0, fourFunc_wire_57_1, fourFunc_wire_57_2});
fanout_n #(3, 0, 0) FANOUT_3 (fourFunc_wire_62, {fourFunc_wire_62_0, fourFunc_wire_62_1, fourFunc_wire_62_2});
fanout_n #(3, 0, 0) FANOUT_4 (fourFunc_wire_67, {fourFunc_wire_67_0, fourFunc_wire_67_1, fourFunc_wire_67_2});
fanout_n #(3, 0, 0) FANOUT_5 (fourFunc_wire_72, {fourFunc_wire_72_0, fourFunc_wire_72_1, fourFunc_wire_72_2});
fanout_n #(3, 0, 0) FANOUT_6 (fourFunc_wire_77, {fourFunc_wire_77_0, fourFunc_wire_77_1, fourFunc_wire_77_2});
fanout_n #(3, 0, 0) FANOUT_7 (fourFunc_wire_87, {fourFunc_wire_87_0, fourFunc_wire_87_1, fourFunc_wire_87_2});
fanout_n #(3, 0, 0) FANOUT_8 (fourFunc_wire_92, {fourFunc_wire_92_0, fourFunc_wire_92_1, fourFunc_wire_92_2});
fanout_n #(3, 0, 0) FANOUT_9 (fourFunc_wire_96, {fourFunc_wire_96_0, fourFunc_wire_96_1, fourFunc_wire_96_2});
fanout_n #(3, 0, 0) FANOUT_10 (fourFunc_wire_100, {fourFunc_wire_100_0, fourFunc_wire_100_1, fourFunc_wire_100_2});
fanout_n #(3, 0, 0) FANOUT_11 (fourFunc_wire_104, {fourFunc_wire_104_0, fourFunc_wire_104_1, fourFunc_wire_104_2});
fanout_n #(3, 0, 0) FANOUT_12 (fourFunc_wire_108, {fourFunc_wire_108_0, fourFunc_wire_108_1, fourFunc_wire_108_2});
fanout_n #(3, 0, 0) FANOUT_13 (fourFunc_wire_116, {fourFunc_wire_116_0, fourFunc_wire_116_1, fourFunc_wire_116_2});
fanout_n #(3, 0, 0) FANOUT_14 (fourFunc_wire_121, {fourFunc_wire_121_0, fourFunc_wire_121_1, fourFunc_wire_121_2});
fanout_n #(3, 0, 0) FANOUT_15 (fourFunc_wire_125, {fourFunc_wire_125_0, fourFunc_wire_125_1, fourFunc_wire_125_2});
fanout_n #(3, 0, 0) FANOUT_16 (fourFunc_wire_129, {fourFunc_wire_129_0, fourFunc_wire_129_1, fourFunc_wire_129_2});
fanout_n #(3, 0, 0) FANOUT_17 (fourFunc_wire_133, {fourFunc_wire_133_0, fourFunc_wire_133_1, fourFunc_wire_133_2});
fanout_n #(3, 0, 0) FANOUT_18 (fourFunc_wire_137, {fourFunc_wire_137_0, fourFunc_wire_137_1, fourFunc_wire_137_2});
fanout_n #(3, 0, 0) FANOUT_19 (fourFunc_wire_145, {fourFunc_wire_145_0, fourFunc_wire_145_1, fourFunc_wire_145_2});
fanout_n #(3, 0, 0) FANOUT_20 (fourFunc_wire_150, {fourFunc_wire_150_0, fourFunc_wire_150_1, fourFunc_wire_150_2});
fanout_n #(3, 0, 0) FANOUT_21 (fourFunc_wire_154, {fourFunc_wire_154_0, fourFunc_wire_154_1, fourFunc_wire_154_2});
fanout_n #(3, 0, 0) FANOUT_22 (fourFunc_wire_158, {fourFunc_wire_158_0, fourFunc_wire_158_1, fourFunc_wire_158_2});
fanout_n #(3, 0, 0) FANOUT_23 (fourFunc_wire_162, {fourFunc_wire_162_0, fourFunc_wire_162_1, fourFunc_wire_162_2});
fanout_n #(3, 0, 0) FANOUT_24 (fourFunc_wire_166, {fourFunc_wire_166_0, fourFunc_wire_166_1, fourFunc_wire_166_2});
fanout_n #(3, 0, 0) FANOUT_25 (fourFunc_wire_174, {fourFunc_wire_174_0, fourFunc_wire_174_1, fourFunc_wire_174_2});
fanout_n #(3, 0, 0) FANOUT_26 (fourFunc_wire_179, {fourFunc_wire_179_0, fourFunc_wire_179_1, fourFunc_wire_179_2});
fanout_n #(3, 0, 0) FANOUT_27 (fourFunc_wire_183, {fourFunc_wire_183_0, fourFunc_wire_183_1, fourFunc_wire_183_2});
fanout_n #(3, 0, 0) FANOUT_28 (fourFunc_wire_187, {fourFunc_wire_187_0, fourFunc_wire_187_1, fourFunc_wire_187_2});
fanout_n #(3, 0, 0) FANOUT_29 (fourFunc_wire_191, {fourFunc_wire_191_0, fourFunc_wire_191_1, fourFunc_wire_191_2});
fanout_n #(3, 0, 0) FANOUT_30 (fourFunc_wire_195, {fourFunc_wire_195_0, fourFunc_wire_195_1, fourFunc_wire_195_2});
fanout_n #(3, 0, 0) FANOUT_31 (fourFunc_wire_203, {fourFunc_wire_203_0, fourFunc_wire_203_1, fourFunc_wire_203_2});
fanout_n #(3, 0, 0) FANOUT_32 (fourFunc_wire_208, {fourFunc_wire_208_0, fourFunc_wire_208_1, fourFunc_wire_208_2});
fanout_n #(3, 0, 0) FANOUT_33 (fourFunc_wire_212, {fourFunc_wire_212_0, fourFunc_wire_212_1, fourFunc_wire_212_2});
fanout_n #(3, 0, 0) FANOUT_34 (fourFunc_wire_216, {fourFunc_wire_216_0, fourFunc_wire_216_1, fourFunc_wire_216_2});
fanout_n #(3, 0, 0) FANOUT_35 (fourFunc_wire_220, {fourFunc_wire_220_0, fourFunc_wire_220_1, fourFunc_wire_220_2});
fanout_n #(3, 0, 0) FANOUT_36 (fourFunc_wire_224, {fourFunc_wire_224_0, fourFunc_wire_224_1, fourFunc_wire_224_2});
fanout_n #(2, 0, 0) FANOUT_37 (fourFunc_wire_84, {fourFunc_wire_84_0, fourFunc_wire_84_1});
fanout_n #(2, 0, 0) FANOUT_38 (fourFunc_wire_79, {fourFunc_wire_79_0, fourFunc_wire_79_1});
fanout_n #(2, 0, 0) FANOUT_39 (fourFunc_wire_74, {fourFunc_wire_74_0, fourFunc_wire_74_1});
fanout_n #(2, 0, 0) FANOUT_40 (fourFunc_wire_69, {fourFunc_wire_69_0, fourFunc_wire_69_1});
fanout_n #(2, 0, 0) FANOUT_41 (fourFunc_wire_64, {fourFunc_wire_64_0, fourFunc_wire_64_1});
fanout_n #(2, 0, 0) FANOUT_42 (fourFunc_wire_59, {fourFunc_wire_59_0, fourFunc_wire_59_1});
fanout_n #(2, 0, 0) FANOUT_43 (fourFunc_wire_56, {fourFunc_wire_56_0, fourFunc_wire_56_1});
fanout_n #(3, 0, 0) FANOUT_44 (fourFunc_wire_91, {fourFunc_wire_91_0, fourFunc_wire_91_1, fourFunc_wire_91_2});
fanout_n #(2, 0, 0) FANOUT_45 (fourFunc_wire_114, {fourFunc_wire_114_0, fourFunc_wire_114_1});
fanout_n #(2, 0, 0) FANOUT_46 (fourFunc_wire_110, {fourFunc_wire_110_0, fourFunc_wire_110_1});
fanout_n #(2, 0, 0) FANOUT_47 (fourFunc_wire_106, {fourFunc_wire_106_0, fourFunc_wire_106_1});
fanout_n #(2, 0, 0) FANOUT_48 (fourFunc_wire_102, {fourFunc_wire_102_0, fourFunc_wire_102_1});
fanout_n #(2, 0, 0) FANOUT_49 (fourFunc_wire_98, {fourFunc_wire_98_0, fourFunc_wire_98_1});
fanout_n #(2, 0, 0) FANOUT_50 (fourFunc_wire_94, {fourFunc_wire_94_0, fourFunc_wire_94_1});
fanout_n #(2, 0, 0) FANOUT_51 (fourFunc_wire_89, {fourFunc_wire_89_0, fourFunc_wire_89_1});
fanout_n #(3, 0, 0) FANOUT_52 (fourFunc_wire_120, {fourFunc_wire_120_0, fourFunc_wire_120_1, fourFunc_wire_120_2});
fanout_n #(2, 0, 0) FANOUT_53 (fourFunc_wire_143, {fourFunc_wire_143_0, fourFunc_wire_143_1});
fanout_n #(2, 0, 0) FANOUT_54 (fourFunc_wire_139, {fourFunc_wire_139_0, fourFunc_wire_139_1});
fanout_n #(2, 0, 0) FANOUT_55 (fourFunc_wire_135, {fourFunc_wire_135_0, fourFunc_wire_135_1});
fanout_n #(2, 0, 0) FANOUT_56 (fourFunc_wire_131, {fourFunc_wire_131_0, fourFunc_wire_131_1});
fanout_n #(2, 0, 0) FANOUT_57 (fourFunc_wire_127, {fourFunc_wire_127_0, fourFunc_wire_127_1});
fanout_n #(2, 0, 0) FANOUT_58 (fourFunc_wire_123, {fourFunc_wire_123_0, fourFunc_wire_123_1});
fanout_n #(2, 0, 0) FANOUT_59 (fourFunc_wire_118, {fourFunc_wire_118_0, fourFunc_wire_118_1});
fanout_n #(3, 0, 0) FANOUT_60 (fourFunc_wire_149, {fourFunc_wire_149_0, fourFunc_wire_149_1, fourFunc_wire_149_2});
fanout_n #(2, 0, 0) FANOUT_61 (fourFunc_wire_172, {fourFunc_wire_172_0, fourFunc_wire_172_1});
fanout_n #(2, 0, 0) FANOUT_62 (fourFunc_wire_168, {fourFunc_wire_168_0, fourFunc_wire_168_1});
fanout_n #(2, 0, 0) FANOUT_63 (fourFunc_wire_164, {fourFunc_wire_164_0, fourFunc_wire_164_1});
fanout_n #(2, 0, 0) FANOUT_64 (fourFunc_wire_160, {fourFunc_wire_160_0, fourFunc_wire_160_1});
fanout_n #(2, 0, 0) FANOUT_65 (fourFunc_wire_156, {fourFunc_wire_156_0, fourFunc_wire_156_1});
fanout_n #(2, 0, 0) FANOUT_66 (fourFunc_wire_152, {fourFunc_wire_152_0, fourFunc_wire_152_1});
fanout_n #(2, 0, 0) FANOUT_67 (fourFunc_wire_147, {fourFunc_wire_147_0, fourFunc_wire_147_1});
fanout_n #(3, 0, 0) FANOUT_68 (fourFunc_wire_178, {fourFunc_wire_178_0, fourFunc_wire_178_1, fourFunc_wire_178_2});
fanout_n #(2, 0, 0) FANOUT_69 (fourFunc_wire_201, {fourFunc_wire_201_0, fourFunc_wire_201_1});
fanout_n #(2, 0, 0) FANOUT_70 (fourFunc_wire_197, {fourFunc_wire_197_0, fourFunc_wire_197_1});
fanout_n #(2, 0, 0) FANOUT_71 (fourFunc_wire_193, {fourFunc_wire_193_0, fourFunc_wire_193_1});
fanout_n #(2, 0, 0) FANOUT_72 (fourFunc_wire_189, {fourFunc_wire_189_0, fourFunc_wire_189_1});
fanout_n #(2, 0, 0) FANOUT_73 (fourFunc_wire_185, {fourFunc_wire_185_0, fourFunc_wire_185_1});
fanout_n #(2, 0, 0) FANOUT_74 (fourFunc_wire_181, {fourFunc_wire_181_0, fourFunc_wire_181_1});
fanout_n #(2, 0, 0) FANOUT_75 (fourFunc_wire_176, {fourFunc_wire_176_0, fourFunc_wire_176_1});
fanout_n #(3, 0, 0) FANOUT_76 (fourFunc_wire_207, {fourFunc_wire_207_0, fourFunc_wire_207_1, fourFunc_wire_207_2});
fanout_n #(2, 0, 0) FANOUT_77 (fourFunc_wire_230, {fourFunc_wire_230_0, fourFunc_wire_230_1});
fanout_n #(2, 0, 0) FANOUT_78 (fourFunc_wire_226, {fourFunc_wire_226_0, fourFunc_wire_226_1});
fanout_n #(2, 0, 0) FANOUT_79 (fourFunc_wire_222, {fourFunc_wire_222_0, fourFunc_wire_222_1});
fanout_n #(2, 0, 0) FANOUT_80 (fourFunc_wire_218, {fourFunc_wire_218_0, fourFunc_wire_218_1});
fanout_n #(2, 0, 0) FANOUT_81 (fourFunc_wire_214, {fourFunc_wire_214_0, fourFunc_wire_214_1});
fanout_n #(2, 0, 0) FANOUT_82 (fourFunc_wire_210, {fourFunc_wire_210_0, fourFunc_wire_210_1});
fanout_n #(2, 0, 0) FANOUT_83 (fourFunc_wire_205, {fourFunc_wire_205_0, fourFunc_wire_205_1});
fanout_n #(3, 0, 0) FANOUT_84 (fourFunc_wire_236, {fourFunc_wire_236_0, fourFunc_wire_236_1, fourFunc_wire_236_2});
fanout_n #(2, 0, 0) FANOUT_85 (fourFunc_wire_259, {fourFunc_wire_259_0, fourFunc_wire_259_1});
fanout_n #(2, 0, 0) FANOUT_86 (fourFunc_wire_255, {fourFunc_wire_255_0, fourFunc_wire_255_1});
fanout_n #(2, 0, 0) FANOUT_87 (fourFunc_wire_251, {fourFunc_wire_251_0, fourFunc_wire_251_1});
fanout_n #(2, 0, 0) FANOUT_88 (fourFunc_wire_247, {fourFunc_wire_247_0, fourFunc_wire_247_1});
fanout_n #(2, 0, 0) FANOUT_89 (fourFunc_wire_243, {fourFunc_wire_243_0, fourFunc_wire_243_1});
fanout_n #(2, 0, 0) FANOUT_90 (fourFunc_wire_239, {fourFunc_wire_239_0, fourFunc_wire_239_1});
fanout_n #(2, 0, 0) FANOUT_91 (fourFunc_wire_234, {fourFunc_wire_234_0, fourFunc_wire_234_1});
fanout_n #(3, 0, 0) FANOUT_92 (fourFunc_wire_61, {fourFunc_wire_61_0, fourFunc_wire_61_1, fourFunc_wire_61_2});
fanout_n #(3, 0, 0) FANOUT_93 (fourFunc_wire_66, {fourFunc_wire_66_0, fourFunc_wire_66_1, fourFunc_wire_66_2});
fanout_n #(3, 0, 0) FANOUT_94 (fourFunc_wire_71, {fourFunc_wire_71_0, fourFunc_wire_71_1, fourFunc_wire_71_2});
fanout_n #(3, 0, 0) FANOUT_95 (fourFunc_wire_76, {fourFunc_wire_76_0, fourFunc_wire_76_1, fourFunc_wire_76_2});
fanout_n #(3, 0, 0) FANOUT_96 (fourFunc_wire_81, {fourFunc_wire_81_0, fourFunc_wire_81_1, fourFunc_wire_81_2});
fanout_n #(3, 0, 0) FANOUT_97 (fourFunc_wire_86, {fourFunc_wire_86_0, fourFunc_wire_86_1, fourFunc_wire_86_2});
fanout_n #(2, 0, 0) FANOUT_98 (fourFunc_wire_261, {fourFunc_wire_261_0, fourFunc_wire_261_1});
fanout_n #(3, 0, 0) FANOUT_99 (fourFunc_wire_60, {fourFunc_wire_60_0, fourFunc_wire_60_1, fourFunc_wire_60_2});
fanout_n #(3, 0, 0) FANOUT_100 (fourFunc_wire_65, {fourFunc_wire_65_0, fourFunc_wire_65_1, fourFunc_wire_65_2});
fanout_n #(3, 0, 0) FANOUT_101 (fourFunc_wire_70, {fourFunc_wire_70_0, fourFunc_wire_70_1, fourFunc_wire_70_2});
fanout_n #(3, 0, 0) FANOUT_102 (fourFunc_wire_75, {fourFunc_wire_75_0, fourFunc_wire_75_1, fourFunc_wire_75_2});
fanout_n #(3, 0, 0) FANOUT_103 (fourFunc_wire_80, {fourFunc_wire_80_0, fourFunc_wire_80_1, fourFunc_wire_80_2});
fanout_n #(3, 0, 0) FANOUT_104 (fourFunc_wire_85, {fourFunc_wire_85_0, fourFunc_wire_85_1, fourFunc_wire_85_2});
fanout_n #(3, 0, 0) FANOUT_105 (fourFunc_wire_90, {fourFunc_wire_90_0, fourFunc_wire_90_1, fourFunc_wire_90_2});
fanout_n #(3, 0, 0) FANOUT_106 (fourFunc_wire_95, {fourFunc_wire_95_0, fourFunc_wire_95_1, fourFunc_wire_95_2});
fanout_n #(3, 0, 0) FANOUT_107 (fourFunc_wire_99, {fourFunc_wire_99_0, fourFunc_wire_99_1, fourFunc_wire_99_2});
fanout_n #(3, 0, 0) FANOUT_108 (fourFunc_wire_103, {fourFunc_wire_103_0, fourFunc_wire_103_1, fourFunc_wire_103_2});
fanout_n #(3, 0, 0) FANOUT_109 (fourFunc_wire_107, {fourFunc_wire_107_0, fourFunc_wire_107_1, fourFunc_wire_107_2});
fanout_n #(3, 0, 0) FANOUT_110 (fourFunc_wire_111, {fourFunc_wire_111_0, fourFunc_wire_111_1, fourFunc_wire_111_2});
fanout_n #(3, 0, 0) FANOUT_111 (fourFunc_wire_115, {fourFunc_wire_115_0, fourFunc_wire_115_1, fourFunc_wire_115_2});
fanout_n #(3, 0, 0) FANOUT_112 (fourFunc_wire_119, {fourFunc_wire_119_0, fourFunc_wire_119_1, fourFunc_wire_119_2});
fanout_n #(3, 0, 0) FANOUT_113 (fourFunc_wire_124, {fourFunc_wire_124_0, fourFunc_wire_124_1, fourFunc_wire_124_2});
fanout_n #(3, 0, 0) FANOUT_114 (fourFunc_wire_128, {fourFunc_wire_128_0, fourFunc_wire_128_1, fourFunc_wire_128_2});
fanout_n #(3, 0, 0) FANOUT_115 (fourFunc_wire_132, {fourFunc_wire_132_0, fourFunc_wire_132_1, fourFunc_wire_132_2});
fanout_n #(3, 0, 0) FANOUT_116 (fourFunc_wire_136, {fourFunc_wire_136_0, fourFunc_wire_136_1, fourFunc_wire_136_2});
fanout_n #(3, 0, 0) FANOUT_117 (fourFunc_wire_140, {fourFunc_wire_140_0, fourFunc_wire_140_1, fourFunc_wire_140_2});
fanout_n #(3, 0, 0) FANOUT_118 (fourFunc_wire_144, {fourFunc_wire_144_0, fourFunc_wire_144_1, fourFunc_wire_144_2});
fanout_n #(3, 0, 0) FANOUT_119 (fourFunc_wire_148, {fourFunc_wire_148_0, fourFunc_wire_148_1, fourFunc_wire_148_2});
fanout_n #(3, 0, 0) FANOUT_120 (fourFunc_wire_153, {fourFunc_wire_153_0, fourFunc_wire_153_1, fourFunc_wire_153_2});
fanout_n #(3, 0, 0) FANOUT_121 (fourFunc_wire_157, {fourFunc_wire_157_0, fourFunc_wire_157_1, fourFunc_wire_157_2});
fanout_n #(3, 0, 0) FANOUT_122 (fourFunc_wire_161, {fourFunc_wire_161_0, fourFunc_wire_161_1, fourFunc_wire_161_2});
fanout_n #(3, 0, 0) FANOUT_123 (fourFunc_wire_165, {fourFunc_wire_165_0, fourFunc_wire_165_1, fourFunc_wire_165_2});
fanout_n #(3, 0, 0) FANOUT_124 (fourFunc_wire_169, {fourFunc_wire_169_0, fourFunc_wire_169_1, fourFunc_wire_169_2});
fanout_n #(3, 0, 0) FANOUT_125 (fourFunc_wire_173, {fourFunc_wire_173_0, fourFunc_wire_173_1, fourFunc_wire_173_2});
fanout_n #(3, 0, 0) FANOUT_126 (fourFunc_wire_177, {fourFunc_wire_177_0, fourFunc_wire_177_1, fourFunc_wire_177_2});
fanout_n #(3, 0, 0) FANOUT_127 (fourFunc_wire_182, {fourFunc_wire_182_0, fourFunc_wire_182_1, fourFunc_wire_182_2});
fanout_n #(3, 0, 0) FANOUT_128 (fourFunc_wire_186, {fourFunc_wire_186_0, fourFunc_wire_186_1, fourFunc_wire_186_2});
fanout_n #(3, 0, 0) FANOUT_129 (fourFunc_wire_190, {fourFunc_wire_190_0, fourFunc_wire_190_1, fourFunc_wire_190_2});
fanout_n #(3, 0, 0) FANOUT_130 (fourFunc_wire_194, {fourFunc_wire_194_0, fourFunc_wire_194_1, fourFunc_wire_194_2});
fanout_n #(3, 0, 0) FANOUT_131 (fourFunc_wire_198, {fourFunc_wire_198_0, fourFunc_wire_198_1, fourFunc_wire_198_2});
fanout_n #(3, 0, 0) FANOUT_132 (fourFunc_wire_202, {fourFunc_wire_202_0, fourFunc_wire_202_1, fourFunc_wire_202_2});
fanout_n #(3, 0, 0) FANOUT_133 (fourFunc_wire_206, {fourFunc_wire_206_0, fourFunc_wire_206_1, fourFunc_wire_206_2});
fanout_n #(3, 0, 0) FANOUT_134 (fourFunc_wire_211, {fourFunc_wire_211_0, fourFunc_wire_211_1, fourFunc_wire_211_2});
fanout_n #(3, 0, 0) FANOUT_135 (fourFunc_wire_215, {fourFunc_wire_215_0, fourFunc_wire_215_1, fourFunc_wire_215_2});
fanout_n #(3, 0, 0) FANOUT_136 (fourFunc_wire_219, {fourFunc_wire_219_0, fourFunc_wire_219_1, fourFunc_wire_219_2});
fanout_n #(3, 0, 0) FANOUT_137 (fourFunc_wire_223, {fourFunc_wire_223_0, fourFunc_wire_223_1, fourFunc_wire_223_2});
fanout_n #(3, 0, 0) FANOUT_138 (fourFunc_wire_227, {fourFunc_wire_227_0, fourFunc_wire_227_1, fourFunc_wire_227_2});
fanout_n #(3, 0, 0) FANOUT_139 (fourFunc_wire_231, {fourFunc_wire_231_0, fourFunc_wire_231_1, fourFunc_wire_231_2});
fanout_n #(3, 0, 0) FANOUT_140 (fourFunc_wire_235, {fourFunc_wire_235_0, fourFunc_wire_235_1, fourFunc_wire_235_2});
fanout_n #(3, 0, 0) FANOUT_141 (fourFunc_wire_240, {fourFunc_wire_240_0, fourFunc_wire_240_1, fourFunc_wire_240_2});
fanout_n #(3, 0, 0) FANOUT_142 (fourFunc_wire_244, {fourFunc_wire_244_0, fourFunc_wire_244_1, fourFunc_wire_244_2});
fanout_n #(3, 0, 0) FANOUT_143 (fourFunc_wire_248, {fourFunc_wire_248_0, fourFunc_wire_248_1, fourFunc_wire_248_2});
fanout_n #(3, 0, 0) FANOUT_144 (fourFunc_wire_252, {fourFunc_wire_252_0, fourFunc_wire_252_1, fourFunc_wire_252_2});
fanout_n #(3, 0, 0) FANOUT_145 (fourFunc_wire_256, {fourFunc_wire_256_0, fourFunc_wire_256_1, fourFunc_wire_256_2});
fanout_n #(3, 0, 0) FANOUT_146 (fourFunc_wire_260, {fourFunc_wire_260_0, fourFunc_wire_260_1, fourFunc_wire_260_2});
fanout_n #(2, 0, 0) FANOUT_147 (fourFunc_wire_502, {fourFunc_wire_502_0, fourFunc_wire_502_1});
fanout_n #(2, 0, 0) FANOUT_148 (fourFunc_wire_499, {fourFunc_wire_499_0, fourFunc_wire_499_1});
fanout_n #(2, 0, 0) FANOUT_149 (fourFunc_wire_496, {fourFunc_wire_496_0, fourFunc_wire_496_1});
fanout_n #(2, 0, 0) FANOUT_150 (fourFunc_wire_493, {fourFunc_wire_493_0, fourFunc_wire_493_1});
fanout_n #(2, 0, 0) FANOUT_151 (fourFunc_wire_490, {fourFunc_wire_490_0, fourFunc_wire_490_1});
fanout_n #(2, 0, 0) FANOUT_152 (fourFunc_wire_487, {fourFunc_wire_487_0, fourFunc_wire_487_1});
fanout_n #(2, 0, 0) FANOUT_153 (fourFunc_wire_484, {fourFunc_wire_484_0, fourFunc_wire_484_1});
fanout_n #(2, 0, 0) FANOUT_154 (fourFunc_wire_479, {fourFunc_wire_479_0, fourFunc_wire_479_1});
fanout_n #(2, 0, 0) FANOUT_155 (fourFunc_wire_475, {fourFunc_wire_475_0, fourFunc_wire_475_1});
fanout_n #(2, 0, 0) FANOUT_156 (fourFunc_wire_471, {fourFunc_wire_471_0, fourFunc_wire_471_1});
fanout_n #(2, 0, 0) FANOUT_157 (fourFunc_wire_467, {fourFunc_wire_467_0, fourFunc_wire_467_1});
fanout_n #(2, 0, 0) FANOUT_158 (fourFunc_wire_463, {fourFunc_wire_463_0, fourFunc_wire_463_1});
fanout_n #(2, 0, 0) FANOUT_159 (fourFunc_wire_459, {fourFunc_wire_459_0, fourFunc_wire_459_1});
fanout_n #(2, 0, 0) FANOUT_160 (fourFunc_wire_455, {fourFunc_wire_455_0, fourFunc_wire_455_1});
fanout_n #(2, 0, 0) FANOUT_161 (fourFunc_wire_451, {fourFunc_wire_451_0, fourFunc_wire_451_1});
fanout_n #(3, 0, 0) FANOUT_162 (fourFunc_wire_448, {fourFunc_wire_448_0, fourFunc_wire_448_1, fourFunc_wire_448_2});
fanout_n #(22, 0, 0) FANOUT_163 (fourFunc_wire_563, {fourFunc_wire_563_0, fourFunc_wire_563_1, fourFunc_wire_563_2, fourFunc_wire_563_3, fourFunc_wire_563_4, fourFunc_wire_563_5, fourFunc_wire_563_6, fourFunc_wire_563_7, fourFunc_wire_563_8, fourFunc_wire_563_9, fourFunc_wire_563_10, fourFunc_wire_563_11, fourFunc_wire_563_12, fourFunc_wire_563_13, fourFunc_wire_563_14, fourFunc_wire_563_15, fourFunc_wire_563_16, fourFunc_wire_563_17, fourFunc_wire_563_18, fourFunc_wire_563_19, fourFunc_wire_563_20, fourFunc_wire_563_21});
fanout_n #(14, 0, 0) FANOUT_164 (fourFunc_wire_11, {fourFunc_wire_11_0, fourFunc_wire_11_1, fourFunc_wire_11_2, fourFunc_wire_11_3, fourFunc_wire_11_4, fourFunc_wire_11_5, fourFunc_wire_11_6, fourFunc_wire_11_7, fourFunc_wire_11_8, fourFunc_wire_11_9, fourFunc_wire_11_10, fourFunc_wire_11_11, fourFunc_wire_11_12, fourFunc_wire_11_13});
fanout_n #(14, 0, 0) FANOUT_165 (fourFunc_wire_3, {fourFunc_wire_3_0, fourFunc_wire_3_1, fourFunc_wire_3_2, fourFunc_wire_3_3, fourFunc_wire_3_4, fourFunc_wire_3_5, fourFunc_wire_3_6, fourFunc_wire_3_7, fourFunc_wire_3_8, fourFunc_wire_3_9, fourFunc_wire_3_10, fourFunc_wire_3_11, fourFunc_wire_3_12, fourFunc_wire_3_13});
fanout_n #(19, 0, 0) FANOUT_166 (fourFunc_wire_2, {fourFunc_wire_2_0, fourFunc_wire_2_1, fourFunc_wire_2_2, fourFunc_wire_2_3, fourFunc_wire_2_4, fourFunc_wire_2_5, fourFunc_wire_2_6, fourFunc_wire_2_7, fourFunc_wire_2_8, fourFunc_wire_2_9, fourFunc_wire_2_10, fourFunc_wire_2_11, fourFunc_wire_2_12, fourFunc_wire_2_13, fourFunc_wire_2_14, fourFunc_wire_2_15, fourFunc_wire_2_16, fourFunc_wire_2_17, fourFunc_wire_2_18});
fanout_n #(2, 0, 0) FANOUT_167 (fourFunc_wire_564, {fourFunc_wire_564_0, fourFunc_wire_564_1});
fanout_n #(2, 0, 0) FANOUT_168 (fourFunc_wire_565, {fourFunc_wire_565_0, fourFunc_wire_565_1});
fanout_n #(2, 0, 0) FANOUT_169 (fourFunc_wire_566, {fourFunc_wire_566_0, fourFunc_wire_566_1});
fanout_n #(2, 0, 0) FANOUT_170 (fourFunc_wire_567, {fourFunc_wire_567_0, fourFunc_wire_567_1});
fanout_n #(2, 0, 0) FANOUT_171 (fourFunc_wire_568, {fourFunc_wire_568_0, fourFunc_wire_568_1});
fanout_n #(2, 0, 0) FANOUT_172 (fourFunc_wire_569, {fourFunc_wire_569_0, fourFunc_wire_569_1});
fanout_n #(2, 0, 0) FANOUT_173 (fourFunc_wire_570, {fourFunc_wire_570_0, fourFunc_wire_570_1});
fanout_n #(2, 0, 0) FANOUT_174 (fourFunc_wire_571, {fourFunc_wire_571_0, fourFunc_wire_571_1});
fanout_n #(12, 0, 0) FANOUT_175 (fourFunc_wire_422, {fourFunc_wire_422_0, fourFunc_wire_422_1, fourFunc_wire_422_2, fourFunc_wire_422_3, fourFunc_wire_422_4, fourFunc_wire_422_5, fourFunc_wire_422_6, fourFunc_wire_422_7, fourFunc_wire_422_8, fourFunc_wire_422_9, fourFunc_wire_422_10, fourFunc_wire_422_11});
fanout_n #(15, 0, 0) FANOUT_176 (fourFunc_wire_430, {fourFunc_wire_430_0, fourFunc_wire_430_1, fourFunc_wire_430_2, fourFunc_wire_430_3, fourFunc_wire_430_4, fourFunc_wire_430_5, fourFunc_wire_430_6, fourFunc_wire_430_7, fourFunc_wire_430_8, fourFunc_wire_430_9, fourFunc_wire_430_10, fourFunc_wire_430_11, fourFunc_wire_430_12, fourFunc_wire_430_13, fourFunc_wire_430_14});
fanout_n #(15, 0, 0) FANOUT_177 (fourFunc_wire_432, {fourFunc_wire_432_0, fourFunc_wire_432_1, fourFunc_wire_432_2, fourFunc_wire_432_3, fourFunc_wire_432_4, fourFunc_wire_432_5, fourFunc_wire_432_6, fourFunc_wire_432_7, fourFunc_wire_432_8, fourFunc_wire_432_9, fourFunc_wire_432_10, fourFunc_wire_432_11, fourFunc_wire_432_12, fourFunc_wire_432_13, fourFunc_wire_432_14});
fanout_n #(15, 0, 0) FANOUT_178 (fourFunc_wire_433, {fourFunc_wire_433_0, fourFunc_wire_433_1, fourFunc_wire_433_2, fourFunc_wire_433_3, fourFunc_wire_433_4, fourFunc_wire_433_5, fourFunc_wire_433_6, fourFunc_wire_433_7, fourFunc_wire_433_8, fourFunc_wire_433_9, fourFunc_wire_433_10, fourFunc_wire_433_11, fourFunc_wire_433_12, fourFunc_wire_433_13, fourFunc_wire_433_14});
fanout_n #(15, 0, 0) FANOUT_179 (fourFunc_wire_434, {fourFunc_wire_434_0, fourFunc_wire_434_1, fourFunc_wire_434_2, fourFunc_wire_434_3, fourFunc_wire_434_4, fourFunc_wire_434_5, fourFunc_wire_434_6, fourFunc_wire_434_7, fourFunc_wire_434_8, fourFunc_wire_434_9, fourFunc_wire_434_10, fourFunc_wire_434_11, fourFunc_wire_434_12, fourFunc_wire_434_13, fourFunc_wire_434_14});
fanout_n #(15, 0, 0) FANOUT_180 (fourFunc_wire_435, {fourFunc_wire_435_0, fourFunc_wire_435_1, fourFunc_wire_435_2, fourFunc_wire_435_3, fourFunc_wire_435_4, fourFunc_wire_435_5, fourFunc_wire_435_6, fourFunc_wire_435_7, fourFunc_wire_435_8, fourFunc_wire_435_9, fourFunc_wire_435_10, fourFunc_wire_435_11, fourFunc_wire_435_12, fourFunc_wire_435_13, fourFunc_wire_435_14});
fanout_n #(15, 0, 0) FANOUT_181 (fourFunc_wire_436, {fourFunc_wire_436_0, fourFunc_wire_436_1, fourFunc_wire_436_2, fourFunc_wire_436_3, fourFunc_wire_436_4, fourFunc_wire_436_5, fourFunc_wire_436_6, fourFunc_wire_436_7, fourFunc_wire_436_8, fourFunc_wire_436_9, fourFunc_wire_436_10, fourFunc_wire_436_11, fourFunc_wire_436_12, fourFunc_wire_436_13, fourFunc_wire_436_14});
fanout_n #(15, 0, 0) FANOUT_182 (fourFunc_wire_437, {fourFunc_wire_437_0, fourFunc_wire_437_1, fourFunc_wire_437_2, fourFunc_wire_437_3, fourFunc_wire_437_4, fourFunc_wire_437_5, fourFunc_wire_437_6, fourFunc_wire_437_7, fourFunc_wire_437_8, fourFunc_wire_437_9, fourFunc_wire_437_10, fourFunc_wire_437_11, fourFunc_wire_437_12, fourFunc_wire_437_13, fourFunc_wire_437_14});
fanout_n #(6, 0, 0) FANOUT_183 (fourFunc_wire_442, {fourFunc_wire_442_0, fourFunc_wire_442_1, fourFunc_wire_442_2, fourFunc_wire_442_3, fourFunc_wire_442_4, fourFunc_wire_442_5});
fanout_n #(8, 0, 0) FANOUT_184 (fourFunc_wire_476, {fourFunc_wire_476_0, fourFunc_wire_476_1, fourFunc_wire_476_2, fourFunc_wire_476_3, fourFunc_wire_476_4, fourFunc_wire_476_5, fourFunc_wire_476_6, fourFunc_wire_476_7});
fanout_n #(8, 0, 0) FANOUT_185 (fourFunc_wire_472, {fourFunc_wire_472_0, fourFunc_wire_472_1, fourFunc_wire_472_2, fourFunc_wire_472_3, fourFunc_wire_472_4, fourFunc_wire_472_5, fourFunc_wire_472_6, fourFunc_wire_472_7});
fanout_n #(8, 0, 0) FANOUT_186 (fourFunc_wire_468, {fourFunc_wire_468_0, fourFunc_wire_468_1, fourFunc_wire_468_2, fourFunc_wire_468_3, fourFunc_wire_468_4, fourFunc_wire_468_5, fourFunc_wire_468_6, fourFunc_wire_468_7});
fanout_n #(8, 0, 0) FANOUT_187 (fourFunc_wire_464, {fourFunc_wire_464_0, fourFunc_wire_464_1, fourFunc_wire_464_2, fourFunc_wire_464_3, fourFunc_wire_464_4, fourFunc_wire_464_5, fourFunc_wire_464_6, fourFunc_wire_464_7});
fanout_n #(8, 0, 0) FANOUT_188 (fourFunc_wire_460, {fourFunc_wire_460_0, fourFunc_wire_460_1, fourFunc_wire_460_2, fourFunc_wire_460_3, fourFunc_wire_460_4, fourFunc_wire_460_5, fourFunc_wire_460_6, fourFunc_wire_460_7});
fanout_n #(8, 0, 0) FANOUT_189 (fourFunc_wire_456, {fourFunc_wire_456_0, fourFunc_wire_456_1, fourFunc_wire_456_2, fourFunc_wire_456_3, fourFunc_wire_456_4, fourFunc_wire_456_5, fourFunc_wire_456_6, fourFunc_wire_456_7});
fanout_n #(8, 0, 0) FANOUT_190 (fourFunc_wire_452, {fourFunc_wire_452_0, fourFunc_wire_452_1, fourFunc_wire_452_2, fourFunc_wire_452_3, fourFunc_wire_452_4, fourFunc_wire_452_5, fourFunc_wire_452_6, fourFunc_wire_452_7});
fanout_n #(7, 0, 0) FANOUT_191 (fourFunc_wire_447, {fourFunc_wire_447_0, fourFunc_wire_447_1, fourFunc_wire_447_2, fourFunc_wire_447_3, fourFunc_wire_447_4, fourFunc_wire_447_5, fourFunc_wire_447_6});
fanout_n #(4, 0, 0) FANOUT_192 (fourFunc_wire_444, {fourFunc_wire_444_0, fourFunc_wire_444_1, fourFunc_wire_444_2, fourFunc_wire_444_3});
fanout_n #(2, 0, 0) FANOUT_193 (fourFunc_wire_594, {fourFunc_wire_594_0, fourFunc_wire_594_1});
fanout_n #(4, 0, 0) FANOUT_194 (fourFunc_wire_600, {fourFunc_wire_600_0, fourFunc_wire_600_1, fourFunc_wire_600_2, fourFunc_wire_600_3});
fanout_n #(5, 0, 0) FANOUT_195 (fourFunc_wire_601, {fourFunc_wire_601_0, fourFunc_wire_601_1, fourFunc_wire_601_2, fourFunc_wire_601_3, fourFunc_wire_601_4});
fanout_n #(3, 0, 0) FANOUT_196 (fourFunc_wire_602, {fourFunc_wire_602_0, fourFunc_wire_602_1, fourFunc_wire_602_2});
fanout_n #(20, 0, 0) FANOUT_197 (fourFunc_wire_598, {fourFunc_wire_598_0, fourFunc_wire_598_1, fourFunc_wire_598_2, fourFunc_wire_598_3, fourFunc_wire_598_4, fourFunc_wire_598_5, fourFunc_wire_598_6, fourFunc_wire_598_7, fourFunc_wire_598_8, fourFunc_wire_598_9, fourFunc_wire_598_10, fourFunc_wire_598_11, fourFunc_wire_598_12, fourFunc_wire_598_13, fourFunc_wire_598_14, fourFunc_wire_598_15, fourFunc_wire_598_16, fourFunc_wire_598_17, fourFunc_wire_598_18, fourFunc_wire_598_19});
fanout_n #(5, 0, 0) FANOUT_198 (fourFunc_wire_593, {fourFunc_wire_593_0, fourFunc_wire_593_1, fourFunc_wire_593_2, fourFunc_wire_593_3, fourFunc_wire_593_4});
fanout_n #(32, 0, 0) FANOUT_199 (fourFunc_wire_611, {fourFunc_wire_611_0, fourFunc_wire_611_1, fourFunc_wire_611_2, fourFunc_wire_611_3, fourFunc_wire_611_4, fourFunc_wire_611_5, fourFunc_wire_611_6, fourFunc_wire_611_7, fourFunc_wire_611_8, fourFunc_wire_611_9, fourFunc_wire_611_10, fourFunc_wire_611_11, fourFunc_wire_611_12, fourFunc_wire_611_13, fourFunc_wire_611_14, fourFunc_wire_611_15, fourFunc_wire_611_16, fourFunc_wire_611_17, fourFunc_wire_611_18, fourFunc_wire_611_19, fourFunc_wire_611_20, fourFunc_wire_611_21, fourFunc_wire_611_22, fourFunc_wire_611_23, fourFunc_wire_611_24, fourFunc_wire_611_25, fourFunc_wire_611_26, fourFunc_wire_611_27, fourFunc_wire_611_28, fourFunc_wire_611_29, fourFunc_wire_611_30, fourFunc_wire_611_31});
fanout_n #(2, 0, 0) FANOUT_200 (fourFunc_wire_612, {fourFunc_wire_612_0, fourFunc_wire_612_1});
fanout_n #(2, 0, 0) FANOUT_201 (fourFunc_wire_618, {fourFunc_wire_618_0, fourFunc_wire_618_1});
fanout_n #(3, 0, 0) FANOUT_202 (fourFunc_wire_622, {fourFunc_wire_622_0, fourFunc_wire_622_1, fourFunc_wire_622_2});
fanout_n #(12, 0, 0) FANOUT_203 (fourFunc_wire_621, {fourFunc_wire_621_0, fourFunc_wire_621_1, fourFunc_wire_621_2, fourFunc_wire_621_3, fourFunc_wire_621_4, fourFunc_wire_621_5, fourFunc_wire_621_6, fourFunc_wire_621_7, fourFunc_wire_621_8, fourFunc_wire_621_9, fourFunc_wire_621_10, fourFunc_wire_621_11});
fanout_n #(40, 0, 0) FANOUT_204 (fourFunc_wire_617, {fourFunc_wire_617_0, fourFunc_wire_617_1, fourFunc_wire_617_2, fourFunc_wire_617_3, fourFunc_wire_617_4, fourFunc_wire_617_5, fourFunc_wire_617_6, fourFunc_wire_617_7, fourFunc_wire_617_8, fourFunc_wire_617_9, fourFunc_wire_617_10, fourFunc_wire_617_11, fourFunc_wire_617_12, fourFunc_wire_617_13, fourFunc_wire_617_14, fourFunc_wire_617_15, fourFunc_wire_617_16, fourFunc_wire_617_17, fourFunc_wire_617_18, fourFunc_wire_617_19, fourFunc_wire_617_20, fourFunc_wire_617_21, fourFunc_wire_617_22, fourFunc_wire_617_23, fourFunc_wire_617_24, fourFunc_wire_617_25, fourFunc_wire_617_26, fourFunc_wire_617_27, fourFunc_wire_617_28, fourFunc_wire_617_29, fourFunc_wire_617_30, fourFunc_wire_617_31, fourFunc_wire_617_32, fourFunc_wire_617_33, fourFunc_wire_617_34, fourFunc_wire_617_35, fourFunc_wire_617_36, fourFunc_wire_617_37, fourFunc_wire_617_38, fourFunc_wire_617_39});
fanout_n #(11, 0, 0) FANOUT_205 (fourFunc_wire_659, {fourFunc_wire_659_0, fourFunc_wire_659_1, fourFunc_wire_659_2, fourFunc_wire_659_3, fourFunc_wire_659_4, fourFunc_wire_659_5, fourFunc_wire_659_6, fourFunc_wire_659_7, fourFunc_wire_659_8, fourFunc_wire_659_9, fourFunc_wire_659_10});
fanout_n #(7, 0, 0) FANOUT_206 (fourFunc_wire_431, {fourFunc_wire_431_0, fourFunc_wire_431_1, fourFunc_wire_431_2, fourFunc_wire_431_3, fourFunc_wire_431_4, fourFunc_wire_431_5, fourFunc_wire_431_6});
fanout_n #(8, 0, 0) FANOUT_207 (fourFunc_wire_429, {fourFunc_wire_429_0, fourFunc_wire_429_1, fourFunc_wire_429_2, fourFunc_wire_429_3, fourFunc_wire_429_4, fourFunc_wire_429_5, fourFunc_wire_429_6, fourFunc_wire_429_7});
fanout_n #(8, 0, 0) FANOUT_208 (fourFunc_wire_428, {fourFunc_wire_428_0, fourFunc_wire_428_1, fourFunc_wire_428_2, fourFunc_wire_428_3, fourFunc_wire_428_4, fourFunc_wire_428_5, fourFunc_wire_428_6, fourFunc_wire_428_7});
fanout_n #(8, 0, 0) FANOUT_209 (fourFunc_wire_427, {fourFunc_wire_427_0, fourFunc_wire_427_1, fourFunc_wire_427_2, fourFunc_wire_427_3, fourFunc_wire_427_4, fourFunc_wire_427_5, fourFunc_wire_427_6, fourFunc_wire_427_7});
fanout_n #(8, 0, 0) FANOUT_210 (fourFunc_wire_426, {fourFunc_wire_426_0, fourFunc_wire_426_1, fourFunc_wire_426_2, fourFunc_wire_426_3, fourFunc_wire_426_4, fourFunc_wire_426_5, fourFunc_wire_426_6, fourFunc_wire_426_7});
fanout_n #(8, 0, 0) FANOUT_211 (fourFunc_wire_425, {fourFunc_wire_425_0, fourFunc_wire_425_1, fourFunc_wire_425_2, fourFunc_wire_425_3, fourFunc_wire_425_4, fourFunc_wire_425_5, fourFunc_wire_425_6, fourFunc_wire_425_7});
fanout_n #(8, 0, 0) FANOUT_212 (fourFunc_wire_424, {fourFunc_wire_424_0, fourFunc_wire_424_1, fourFunc_wire_424_2, fourFunc_wire_424_3, fourFunc_wire_424_4, fourFunc_wire_424_5, fourFunc_wire_424_6, fourFunc_wire_424_7});
fanout_n #(8, 0, 0) FANOUT_213 (fourFunc_wire_423, {fourFunc_wire_423_0, fourFunc_wire_423_1, fourFunc_wire_423_2, fourFunc_wire_423_3, fourFunc_wire_423_4, fourFunc_wire_423_5, fourFunc_wire_423_6, fourFunc_wire_423_7});
fanout_n #(9, 0, 0) FANOUT_214 (fourFunc_wire_733, {fourFunc_wire_733_0, fourFunc_wire_733_1, fourFunc_wire_733_2, fourFunc_wire_733_3, fourFunc_wire_733_4, fourFunc_wire_733_5, fourFunc_wire_733_6, fourFunc_wire_733_7, fourFunc_wire_733_8});
fanout_n #(32, 0, 0) FANOUT_215 (fourFunc_wire_7, {fourFunc_wire_7_0, fourFunc_wire_7_1, fourFunc_wire_7_2, fourFunc_wire_7_3, fourFunc_wire_7_4, fourFunc_wire_7_5, fourFunc_wire_7_6, fourFunc_wire_7_7, fourFunc_wire_7_8, fourFunc_wire_7_9, fourFunc_wire_7_10, fourFunc_wire_7_11, fourFunc_wire_7_12, fourFunc_wire_7_13, fourFunc_wire_7_14, fourFunc_wire_7_15, fourFunc_wire_7_16, fourFunc_wire_7_17, fourFunc_wire_7_18, fourFunc_wire_7_19, fourFunc_wire_7_20, fourFunc_wire_7_21, fourFunc_wire_7_22, fourFunc_wire_7_23, fourFunc_wire_7_24, fourFunc_wire_7_25, fourFunc_wire_7_26, fourFunc_wire_7_27, fourFunc_wire_7_28, fourFunc_wire_7_29, fourFunc_wire_7_30, fourFunc_wire_7_31});
fanout_n #(6, 0, 0) FANOUT_216 (fourFunc_wire_610, {fourFunc_wire_610_0, fourFunc_wire_610_1, fourFunc_wire_610_2, fourFunc_wire_610_3, fourFunc_wire_610_4, fourFunc_wire_610_5});
fanout_n #(3, 0, 0) FANOUT_217 (fourFunc_wire_650, {fourFunc_wire_650_0, fourFunc_wire_650_1, fourFunc_wire_650_2});
fanout_n #(3, 0, 0) FANOUT_218 (fourFunc_wire_637, {fourFunc_wire_637_0, fourFunc_wire_637_1, fourFunc_wire_637_2});
fanout_n #(3, 0, 0) FANOUT_219 (fourFunc_wire_639, {fourFunc_wire_639_0, fourFunc_wire_639_1, fourFunc_wire_639_2});
fanout_n #(3, 0, 0) FANOUT_220 (fourFunc_wire_641, {fourFunc_wire_641_0, fourFunc_wire_641_1, fourFunc_wire_641_2});
fanout_n #(3, 0, 0) FANOUT_221 (fourFunc_wire_635, {fourFunc_wire_635_0, fourFunc_wire_635_1, fourFunc_wire_635_2});
fanout_n #(3, 0, 0) FANOUT_222 (fourFunc_wire_643, {fourFunc_wire_643_0, fourFunc_wire_643_1, fourFunc_wire_643_2});
fanout_n #(3, 0, 0) FANOUT_223 (fourFunc_wire_645, {fourFunc_wire_645_0, fourFunc_wire_645_1, fourFunc_wire_645_2});
fanout_n #(3, 0, 0) FANOUT_224 (fourFunc_wire_647, {fourFunc_wire_647_0, fourFunc_wire_647_1, fourFunc_wire_647_2});
fanout_n #(3, 0, 0) FANOUT_225 (fourFunc_wire_649, {fourFunc_wire_649_0, fourFunc_wire_649_1, fourFunc_wire_649_2});
fanout_n #(2, 0, 0) FANOUT_226 (NOT_intermediateXXXwire_735, {NOT_intermediateXXXwire_735_0, NOT_intermediateXXXwire_735_1});
fanout_n #(8, 0, 0) FANOUT_227 (NOT_intermediateXXXwire_739, {NOT_intermediateXXXwire_739_0, NOT_intermediateXXXwire_739_1, NOT_intermediateXXXwire_739_2, NOT_intermediateXXXwire_739_3, NOT_intermediateXXXwire_739_4, NOT_intermediateXXXwire_739_5, NOT_intermediateXXXwire_739_6, NOT_intermediateXXXwire_739_7});
fanout_n #(8, 0, 0) FANOUT_228 (NOT_intermediateXXXwire_963, {NOT_intermediateXXXwire_963_0, NOT_intermediateXXXwire_963_1, NOT_intermediateXXXwire_963_2, NOT_intermediateXXXwire_963_3, NOT_intermediateXXXwire_963_4, NOT_intermediateXXXwire_963_5, NOT_intermediateXXXwire_963_6, NOT_intermediateXXXwire_963_7});
fanout_n #(10, 0, 0) FANOUT_229 (NOT_intermediateXXXwire_834, {NOT_intermediateXXXwire_834_0, NOT_intermediateXXXwire_834_1, NOT_intermediateXXXwire_834_2, NOT_intermediateXXXwire_834_3, NOT_intermediateXXXwire_834_4, NOT_intermediateXXXwire_834_5, NOT_intermediateXXXwire_834_6, NOT_intermediateXXXwire_834_7, NOT_intermediateXXXwire_834_8, NOT_intermediateXXXwire_834_9});


and_n #(2, 0, 0) AND_1 (fourFunc_wire_1, {fourFunc_wire_2_0, fourFunc_wire_3_0});
or_n #(2, 0, 0) OR_1 (fourFunc_wire_4, {fourFunc_wire_1, fourFunc_wire_5});
and_n #(2, 0, 0) AND_2 (fourFunc_wire_6, {fourFunc_wire_2_1, fourFunc_wire_7_0});
or_n #(2, 0, 0) OR_2 (fourFunc_wire_8, {fourFunc_wire_6, fourFunc_wire_9});
nor_n #(2, 0, 0) NOR_1 (fourFunc_wire_9, {fourFunc_wire_2_2, fourFunc_wire_7_1});
notg #(0, 0) NOT_1 (fourFunc_wire_10, fourFunc_wire_11_0);
and_n #(2, 0, 0) AND_3 (fourFunc_wire_5, {fourFunc_wire_10, fourFunc_wire_8});
notg #(0, 0) NOT_2 (fourFunc_wire_12, fourFunc_wire_2_3);
and_n #(2, 0, 0) AND_4 (fourFunc_wire_13, {fourFunc_wire_12, fourFunc_wire_3_1});
nor_n #(2, 0, 0) NOR_2 (fourFunc_wire_14, {fourFunc_wire_3_2, fourFunc_wire_7_2});
nor_n #(2, 0, 0) NOR_3 (fourFunc_wire_15, {fourFunc_wire_2_4, fourFunc_wire_7_3});
or_n #(2, 0, 0) OR_3 (fourFunc_wire_16, {fourFunc_wire_13, fourFunc_wire_14});
or_n #(2, 0, 0) OR_4 (fourFunc_wire_17, {fourFunc_wire_15, fourFunc_wire_18});
and_n #(2, 0, 0) AND_5 (fourFunc_wire_18, {fourFunc_wire_16, fourFunc_wire_11_1});
notg #(0, 0) NOT_3 (fourFunc_wire_19, fourFunc_wire_7_4);
or_n #(2, 0, 0) OR_5 (fourFunc_wire_20, {fourFunc_wire_19, fourFunc_wire_2_5});
notg #(0, 0) NOT_4 (fourFunc_wire_21, fourFunc_wire_3_3);
and_n #(2, 0, 0) AND_6 (fourFunc_wire_22, {fourFunc_wire_21, fourFunc_wire_20});
or_n #(2, 0, 0) OR_6 (fourFunc_wire_23, {fourFunc_wire_22, fourFunc_wire_24});
and_n #(2, 0, 0) AND_7 (fourFunc_wire_25, {fourFunc_wire_23, fourFunc_wire_26});
or_n #(2, 0, 0) OR_7 (fourFunc_wire_27, {fourFunc_wire_25, fourFunc_wire_28});
and_n #(2, 0, 0) AND_8 (fourFunc_wire_29, {fourFunc_wire_3_4, fourFunc_wire_7_5});
and_n #(2, 0, 0) AND_9 (fourFunc_wire_24, {fourFunc_wire_29, fourFunc_wire_30});
notg #(0, 0) NOT_5 (fourFunc_wire_30, fourFunc_wire_2_6);
notg #(0, 0) NOT_6 (fourFunc_wire_26, fourFunc_wire_11_2);
notg #(0, 0) NOT_7 (fourFunc_wire_31, fourFunc_wire_3_5);
and_n #(3, 0, 0) AND_10 (fourFunc_wire_28, {fourFunc_wire_31, fourFunc_wire_32, fourFunc_wire_2_7});
notg #(0, 0) NOT_8 (fourFunc_wire_32, fourFunc_wire_7_6);
nand_n #(2, 0, 0) NAND_1 (fourFunc_wire_33, {fourFunc_wire_11_3, fourFunc_wire_2_8});
notg #(0, 0) NOT_9 (fourFunc_wire_34, fourFunc_wire_7_7);
and_n #(2, 0, 0) AND_11 (fourFunc_wire_35, {fourFunc_wire_34, fourFunc_wire_33});
and_n #(3, 0, 0) AND_12 (fourFunc_wire_36, {fourFunc_wire_11_4, fourFunc_wire_2_9, fourFunc_wire_7_8});
or_n #(2, 0, 0) OR_8 (fourFunc_wire_37, {fourFunc_wire_36, fourFunc_wire_35});
notg #(0, 0) NOT_10 (fourFunc_wire_38, fourFunc_wire_3_6);
and_n #(2, 0, 0) AND_13 (fourFunc_wire_39, {fourFunc_wire_38, fourFunc_wire_37});
and_n #(2, 0, 0) AND_14 (fourFunc_wire_40, {fourFunc_wire_2_10, fourFunc_wire_7_9});
or_n #(2, 0, 0) OR_9 (fourFunc_wire_41, {fourFunc_wire_40, fourFunc_wire_42});
nor_n #(2, 0, 0) NOR_4 (fourFunc_wire_42, {fourFunc_wire_2_11, fourFunc_wire_7_10});
notg #(0, 0) NOT_11 (fourFunc_wire_43, fourFunc_wire_3_7);
and_n #(3, 0, 0) AND_15 (fourFunc_wire_44, {fourFunc_wire_43, fourFunc_wire_45, fourFunc_wire_41});
notg #(0, 0) NOT_12 (fourFunc_wire_45, fourFunc_wire_11_5);
nor_n #(3, 0, 0) NOR_5 (fourFunc_wire_46, {fourFunc_wire_3_8, fourFunc_wire_2_12, fourFunc_wire_7_11});
and_n #(2, 0, 0) AND_16 (fourFunc_wire_47, {fourFunc_wire_11_6, fourFunc_wire_7_12});
or_n #(2, 0, 0) OR_10 (fourFunc_wire_48, {fourFunc_wire_47, fourFunc_wire_49});
nor_n #(2, 0, 0) NOR_6 (fourFunc_wire_49, {fourFunc_wire_11_7, fourFunc_wire_7_13});
notg #(0, 0) NOT_13 (fourFunc_wire_50, fourFunc_wire_3_9);
and_n #(3, 0, 0) AND_17 (fourFunc_wire_51, {fourFunc_wire_50, fourFunc_wire_52, fourFunc_wire_48});
notg #(0, 0) NOT_14 (fourFunc_wire_52, fourFunc_wire_2_13);
nor_n #(4, 0, 0) NOR_7 (fourFunc_wire_53, {fourFunc_wire_11_8, fourFunc_wire_2_14, fourFunc_wire_3_10, fourFunc_wire_7_14});
xor_n #(2, 0, 0) XOR_1 (fourFunc_wire_54, {fourFunc_wire_55, fourFunc_wire_56_0});
xor_n #(2, 0, 0) XOR_2 (fourFunc_wire_57, {fourFunc_wire_58, fourFunc_wire_59_0});
xor_n #(2, 0, 0) XOR_3 (fourFunc_wire_58, {fourFunc_wire_60_0, fourFunc_wire_61_0});
xor_n #(2, 0, 0) XOR_4 (fourFunc_wire_62, {fourFunc_wire_63, fourFunc_wire_64_0});
xor_n #(2, 0, 0) XOR_5 (fourFunc_wire_63, {fourFunc_wire_65_0, fourFunc_wire_66_0});
xor_n #(2, 0, 0) XOR_6 (fourFunc_wire_67, {fourFunc_wire_68, fourFunc_wire_69_0});
xor_n #(2, 0, 0) XOR_7 (fourFunc_wire_68, {fourFunc_wire_70_0, fourFunc_wire_71_0});
xor_n #(2, 0, 0) XOR_8 (fourFunc_wire_72, {fourFunc_wire_73, fourFunc_wire_74_0});
xor_n #(2, 0, 0) XOR_9 (fourFunc_wire_73, {fourFunc_wire_75_0, fourFunc_wire_76_0});
xor_n #(2, 0, 0) XOR_10 (fourFunc_wire_77, {fourFunc_wire_78, fourFunc_wire_79_0});
xor_n #(2, 0, 0) XOR_11 (fourFunc_wire_78, {fourFunc_wire_80_0, fourFunc_wire_81_0});
xor_n #(2, 0, 0) XOR_12 (fourFunc_wire_82, {fourFunc_wire_83, fourFunc_wire_84_0});
xor_n #(2, 0, 0) XOR_13 (fourFunc_wire_83, {fourFunc_wire_85_0, fourFunc_wire_86_0});
xor_n #(2, 0, 0) XOR_14 (fourFunc_wire_87, {fourFunc_wire_88, fourFunc_wire_89_0});
xor_n #(2, 0, 0) XOR_15 (fourFunc_wire_88, {fourFunc_wire_90_0, fourFunc_wire_91_0});
xor_n #(2, 0, 0) XOR_16 (fourFunc_wire_92, {fourFunc_wire_93, fourFunc_wire_94_0});
xor_n #(2, 0, 0) XOR_17 (fourFunc_wire_93, {fourFunc_wire_95_0, fourFunc_wire_54_0});
xor_n #(2, 0, 0) XOR_18 (fourFunc_wire_96, {fourFunc_wire_97, fourFunc_wire_98_0});
xor_n #(2, 0, 0) XOR_19 (fourFunc_wire_97, {fourFunc_wire_99_0, fourFunc_wire_57_0});
xor_n #(2, 0, 0) XOR_20 (fourFunc_wire_100, {fourFunc_wire_101, fourFunc_wire_102_0});
xor_n #(2, 0, 0) XOR_21 (fourFunc_wire_101, {fourFunc_wire_103_0, fourFunc_wire_62_0});
xor_n #(2, 0, 0) XOR_22 (fourFunc_wire_104, {fourFunc_wire_105, fourFunc_wire_106_0});
xor_n #(2, 0, 0) XOR_23 (fourFunc_wire_105, {fourFunc_wire_107_0, fourFunc_wire_67_0});
xor_n #(2, 0, 0) XOR_24 (fourFunc_wire_108, {fourFunc_wire_109, fourFunc_wire_110_0});
xor_n #(2, 0, 0) XOR_25 (fourFunc_wire_109, {fourFunc_wire_111_0, fourFunc_wire_72_0});
xor_n #(2, 0, 0) XOR_26 (fourFunc_wire_112, {fourFunc_wire_113, fourFunc_wire_114_0});
xor_n #(2, 0, 0) XOR_27 (fourFunc_wire_113, {fourFunc_wire_115_0, fourFunc_wire_77_0});
xor_n #(2, 0, 0) XOR_28 (fourFunc_wire_116, {fourFunc_wire_117, fourFunc_wire_118_0});
xor_n #(2, 0, 0) XOR_29 (fourFunc_wire_117, {fourFunc_wire_119_0, fourFunc_wire_120_0});
xor_n #(2, 0, 0) XOR_30 (fourFunc_wire_121, {fourFunc_wire_122, fourFunc_wire_123_0});
xor_n #(2, 0, 0) XOR_31 (fourFunc_wire_122, {fourFunc_wire_124_0, fourFunc_wire_87_0});
xor_n #(2, 0, 0) XOR_32 (fourFunc_wire_125, {fourFunc_wire_126, fourFunc_wire_127_0});
xor_n #(2, 0, 0) XOR_33 (fourFunc_wire_126, {fourFunc_wire_128_0, fourFunc_wire_92_0});
xor_n #(2, 0, 0) XOR_34 (fourFunc_wire_129, {fourFunc_wire_130, fourFunc_wire_131_0});
xor_n #(2, 0, 0) XOR_35 (fourFunc_wire_130, {fourFunc_wire_132_0, fourFunc_wire_96_0});
xor_n #(2, 0, 0) XOR_36 (fourFunc_wire_133, {fourFunc_wire_134, fourFunc_wire_135_0});
xor_n #(2, 0, 0) XOR_37 (fourFunc_wire_134, {fourFunc_wire_136_0, fourFunc_wire_100_0});
xor_n #(2, 0, 0) XOR_38 (fourFunc_wire_137, {fourFunc_wire_138, fourFunc_wire_139_0});
xor_n #(2, 0, 0) XOR_39 (fourFunc_wire_138, {fourFunc_wire_140_0, fourFunc_wire_104_0});
xor_n #(2, 0, 0) XOR_40 (fourFunc_wire_141, {fourFunc_wire_142, fourFunc_wire_143_0});
xor_n #(2, 0, 0) XOR_41 (fourFunc_wire_142, {fourFunc_wire_144_0, fourFunc_wire_108_0});
xor_n #(2, 0, 0) XOR_42 (fourFunc_wire_145, {fourFunc_wire_146, fourFunc_wire_147_0});
xor_n #(2, 0, 0) XOR_43 (fourFunc_wire_146, {fourFunc_wire_148_0, fourFunc_wire_149_0});
xor_n #(2, 0, 0) XOR_44 (fourFunc_wire_150, {fourFunc_wire_151, fourFunc_wire_152_0});
xor_n #(2, 0, 0) XOR_45 (fourFunc_wire_151, {fourFunc_wire_153_0, fourFunc_wire_116_0});
xor_n #(2, 0, 0) XOR_46 (fourFunc_wire_154, {fourFunc_wire_155, fourFunc_wire_156_0});
xor_n #(2, 0, 0) XOR_47 (fourFunc_wire_155, {fourFunc_wire_157_0, fourFunc_wire_121_0});
xor_n #(2, 0, 0) XOR_48 (fourFunc_wire_158, {fourFunc_wire_159, fourFunc_wire_160_0});
xor_n #(2, 0, 0) XOR_49 (fourFunc_wire_159, {fourFunc_wire_161_0, fourFunc_wire_125_0});
xor_n #(2, 0, 0) XOR_50 (fourFunc_wire_162, {fourFunc_wire_163, fourFunc_wire_164_0});
xor_n #(2, 0, 0) XOR_51 (fourFunc_wire_163, {fourFunc_wire_165_0, fourFunc_wire_129_0});
xor_n #(2, 0, 0) XOR_52 (fourFunc_wire_166, {fourFunc_wire_167, fourFunc_wire_168_0});
xor_n #(2, 0, 0) XOR_53 (fourFunc_wire_167, {fourFunc_wire_169_0, fourFunc_wire_133_0});
xor_n #(2, 0, 0) XOR_54 (fourFunc_wire_170, {fourFunc_wire_171, fourFunc_wire_172_0});
xor_n #(2, 0, 0) XOR_55 (fourFunc_wire_171, {fourFunc_wire_173_0, fourFunc_wire_137_0});
xor_n #(2, 0, 0) XOR_56 (fourFunc_wire_174, {fourFunc_wire_175, fourFunc_wire_176_0});
xor_n #(2, 0, 0) XOR_57 (fourFunc_wire_175, {fourFunc_wire_177_0, fourFunc_wire_178_0});
xor_n #(2, 0, 0) XOR_58 (fourFunc_wire_179, {fourFunc_wire_180, fourFunc_wire_181_0});
xor_n #(2, 0, 0) XOR_59 (fourFunc_wire_180, {fourFunc_wire_182_0, fourFunc_wire_145_0});
xor_n #(2, 0, 0) XOR_60 (fourFunc_wire_183, {fourFunc_wire_184, fourFunc_wire_185_0});
xor_n #(2, 0, 0) XOR_61 (fourFunc_wire_184, {fourFunc_wire_186_0, fourFunc_wire_150_0});
xor_n #(2, 0, 0) XOR_62 (fourFunc_wire_187, {fourFunc_wire_188, fourFunc_wire_189_0});
xor_n #(2, 0, 0) XOR_63 (fourFunc_wire_188, {fourFunc_wire_190_0, fourFunc_wire_154_0});
xor_n #(2, 0, 0) XOR_64 (fourFunc_wire_191, {fourFunc_wire_192, fourFunc_wire_193_0});
xor_n #(2, 0, 0) XOR_65 (fourFunc_wire_192, {fourFunc_wire_194_0, fourFunc_wire_158_0});
xor_n #(2, 0, 0) XOR_66 (fourFunc_wire_195, {fourFunc_wire_196, fourFunc_wire_197_0});
xor_n #(2, 0, 0) XOR_67 (fourFunc_wire_196, {fourFunc_wire_198_0, fourFunc_wire_162_0});
xor_n #(2, 0, 0) XOR_68 (fourFunc_wire_199, {fourFunc_wire_200, fourFunc_wire_201_0});
xor_n #(2, 0, 0) XOR_69 (fourFunc_wire_200, {fourFunc_wire_202_0, fourFunc_wire_166_0});
xor_n #(2, 0, 0) XOR_70 (fourFunc_wire_203, {fourFunc_wire_204, fourFunc_wire_205_0});
xor_n #(2, 0, 0) XOR_71 (fourFunc_wire_204, {fourFunc_wire_206_0, fourFunc_wire_207_0});
xor_n #(2, 0, 0) XOR_72 (fourFunc_wire_208, {fourFunc_wire_209, fourFunc_wire_210_0});
xor_n #(2, 0, 0) XOR_73 (fourFunc_wire_209, {fourFunc_wire_211_0, fourFunc_wire_174_0});
xor_n #(2, 0, 0) XOR_74 (fourFunc_wire_212, {fourFunc_wire_213, fourFunc_wire_214_0});
xor_n #(2, 0, 0) XOR_75 (fourFunc_wire_213, {fourFunc_wire_215_0, fourFunc_wire_179_0});
xor_n #(2, 0, 0) XOR_76 (fourFunc_wire_216, {fourFunc_wire_217, fourFunc_wire_218_0});
xor_n #(2, 0, 0) XOR_77 (fourFunc_wire_217, {fourFunc_wire_219_0, fourFunc_wire_183_0});
xor_n #(2, 0, 0) XOR_78 (fourFunc_wire_220, {fourFunc_wire_221, fourFunc_wire_222_0});
xor_n #(2, 0, 0) XOR_79 (fourFunc_wire_221, {fourFunc_wire_223_0, fourFunc_wire_187_0});
xor_n #(2, 0, 0) XOR_80 (fourFunc_wire_224, {fourFunc_wire_225, fourFunc_wire_226_0});
xor_n #(2, 0, 0) XOR_81 (fourFunc_wire_225, {fourFunc_wire_227_0, fourFunc_wire_191_0});
xor_n #(2, 0, 0) XOR_82 (fourFunc_wire_228, {fourFunc_wire_229, fourFunc_wire_230_0});
xor_n #(2, 0, 0) XOR_83 (fourFunc_wire_229, {fourFunc_wire_231_0, fourFunc_wire_195_0});
xor_n #(2, 0, 0) XOR_84 (fourFunc_wire_232, {fourFunc_wire_233, fourFunc_wire_234_0});
xor_n #(2, 0, 0) XOR_85 (fourFunc_wire_233, {fourFunc_wire_235_0, fourFunc_wire_236_0});
xor_n #(2, 0, 0) XOR_86 (fourFunc_wire_237, {fourFunc_wire_238, fourFunc_wire_239_0});
xor_n #(2, 0, 0) XOR_87 (fourFunc_wire_238, {fourFunc_wire_240_0, fourFunc_wire_203_0});
xor_n #(2, 0, 0) XOR_88 (fourFunc_wire_241, {fourFunc_wire_242, fourFunc_wire_243_0});
xor_n #(2, 0, 0) XOR_89 (fourFunc_wire_242, {fourFunc_wire_244_0, fourFunc_wire_208_0});
xor_n #(2, 0, 0) XOR_90 (fourFunc_wire_245, {fourFunc_wire_246, fourFunc_wire_247_0});
xor_n #(2, 0, 0) XOR_91 (fourFunc_wire_246, {fourFunc_wire_248_0, fourFunc_wire_212_0});
xor_n #(2, 0, 0) XOR_92 (fourFunc_wire_249, {fourFunc_wire_250, fourFunc_wire_251_0});
xor_n #(2, 0, 0) XOR_93 (fourFunc_wire_250, {fourFunc_wire_252_0, fourFunc_wire_216_0});
xor_n #(2, 0, 0) XOR_94 (fourFunc_wire_253, {fourFunc_wire_254, fourFunc_wire_255_0});
xor_n #(2, 0, 0) XOR_95 (fourFunc_wire_254, {fourFunc_wire_256_0, fourFunc_wire_220_0});
xor_n #(2, 0, 0) XOR_96 (fourFunc_wire_257, {fourFunc_wire_258, fourFunc_wire_259_0});
xor_n #(2, 0, 0) XOR_97 (fourFunc_wire_258, {fourFunc_wire_260_0, fourFunc_wire_224_0});
bufg #(0, 0) BUF_1 (fourFunc_wire_55, fourFunc_wire_261_0);
and_n #(2, 0, 0) AND_18 (fourFunc_wire_84, {fourFunc_wire_262, fourFunc_wire_263});
and_n #(2, 0, 0) AND_19 (fourFunc_wire_264, {fourFunc_wire_84_1, fourFunc_wire_265});
or_n #(2, 0, 0) OR_11 (fourFunc_wire_79, {fourFunc_wire_266, fourFunc_wire_264});
and_n #(2, 0, 0) AND_20 (fourFunc_wire_267, {fourFunc_wire_79_1, fourFunc_wire_268});
and_n #(2, 0, 0) AND_21 (fourFunc_wire_266, {fourFunc_wire_86_1, fourFunc_wire_85_1});
or_n #(2, 0, 0) OR_12 (fourFunc_wire_265, {fourFunc_wire_86_2, fourFunc_wire_85_2});
or_n #(2, 0, 0) OR_13 (fourFunc_wire_74, {fourFunc_wire_269, fourFunc_wire_267});
and_n #(2, 0, 0) AND_22 (fourFunc_wire_270, {fourFunc_wire_74_1, fourFunc_wire_271});
and_n #(2, 0, 0) AND_23 (fourFunc_wire_269, {fourFunc_wire_81_1, fourFunc_wire_80_1});
or_n #(2, 0, 0) OR_14 (fourFunc_wire_268, {fourFunc_wire_81_2, fourFunc_wire_80_2});
or_n #(2, 0, 0) OR_15 (fourFunc_wire_69, {fourFunc_wire_272, fourFunc_wire_270});
and_n #(2, 0, 0) AND_24 (fourFunc_wire_273, {fourFunc_wire_69_1, fourFunc_wire_274});
and_n #(2, 0, 0) AND_25 (fourFunc_wire_272, {fourFunc_wire_76_1, fourFunc_wire_75_1});
or_n #(2, 0, 0) OR_16 (fourFunc_wire_271, {fourFunc_wire_76_2, fourFunc_wire_75_2});
or_n #(2, 0, 0) OR_17 (fourFunc_wire_64, {fourFunc_wire_275, fourFunc_wire_273});
and_n #(2, 0, 0) AND_26 (fourFunc_wire_276, {fourFunc_wire_64_1, fourFunc_wire_277});
and_n #(2, 0, 0) AND_27 (fourFunc_wire_275, {fourFunc_wire_71_1, fourFunc_wire_70_1});
or_n #(2, 0, 0) OR_18 (fourFunc_wire_274, {fourFunc_wire_71_2, fourFunc_wire_70_2});
or_n #(2, 0, 0) OR_19 (fourFunc_wire_59, {fourFunc_wire_278, fourFunc_wire_276});
and_n #(2, 0, 0) AND_28 (fourFunc_wire_279, {fourFunc_wire_59_1, fourFunc_wire_280});
and_n #(2, 0, 0) AND_29 (fourFunc_wire_278, {fourFunc_wire_66_1, fourFunc_wire_65_1});
or_n #(2, 0, 0) OR_20 (fourFunc_wire_277, {fourFunc_wire_66_2, fourFunc_wire_65_2});
and_n #(2, 0, 0) AND_30 (fourFunc_wire_281, {fourFunc_wire_56_1, fourFunc_wire_261_1});
or_n #(2, 0, 0) OR_21 (fourFunc_wire_56, {fourFunc_wire_282, fourFunc_wire_279});
and_n #(2, 0, 0) AND_31 (fourFunc_wire_282, {fourFunc_wire_61_1, fourFunc_wire_60_1});
or_n #(2, 0, 0) OR_22 (fourFunc_wire_280, {fourFunc_wire_61_2, fourFunc_wire_60_2});
bufg #(0, 0) BUF_2 (fourFunc_wire_91, fourFunc_wire_281);
and_n #(2, 0, 0) AND_32 (fourFunc_wire_114, {fourFunc_wire_82, fourFunc_wire_283});
and_n #(2, 0, 0) AND_33 (fourFunc_wire_284, {fourFunc_wire_114_1, fourFunc_wire_285});
or_n #(2, 0, 0) OR_23 (fourFunc_wire_110, {fourFunc_wire_286, fourFunc_wire_284});
and_n #(2, 0, 0) AND_34 (fourFunc_wire_287, {fourFunc_wire_110_1, fourFunc_wire_288});
and_n #(2, 0, 0) AND_35 (fourFunc_wire_286, {fourFunc_wire_77_1, fourFunc_wire_115_1});
or_n #(2, 0, 0) OR_24 (fourFunc_wire_285, {fourFunc_wire_77_2, fourFunc_wire_115_2});
or_n #(2, 0, 0) OR_25 (fourFunc_wire_106, {fourFunc_wire_289, fourFunc_wire_287});
and_n #(2, 0, 0) AND_36 (fourFunc_wire_290, {fourFunc_wire_106_1, fourFunc_wire_291});
and_n #(2, 0, 0) AND_37 (fourFunc_wire_289, {fourFunc_wire_72_1, fourFunc_wire_111_1});
or_n #(2, 0, 0) OR_26 (fourFunc_wire_288, {fourFunc_wire_72_2, fourFunc_wire_111_2});
or_n #(2, 0, 0) OR_27 (fourFunc_wire_102, {fourFunc_wire_292, fourFunc_wire_290});
and_n #(2, 0, 0) AND_38 (fourFunc_wire_293, {fourFunc_wire_102_1, fourFunc_wire_294});
and_n #(2, 0, 0) AND_39 (fourFunc_wire_292, {fourFunc_wire_67_1, fourFunc_wire_107_1});
or_n #(2, 0, 0) OR_28 (fourFunc_wire_291, {fourFunc_wire_67_2, fourFunc_wire_107_2});
or_n #(2, 0, 0) OR_29 (fourFunc_wire_98, {fourFunc_wire_295, fourFunc_wire_293});
and_n #(2, 0, 0) AND_40 (fourFunc_wire_296, {fourFunc_wire_98_1, fourFunc_wire_297});
and_n #(2, 0, 0) AND_41 (fourFunc_wire_295, {fourFunc_wire_62_1, fourFunc_wire_103_1});
or_n #(2, 0, 0) OR_30 (fourFunc_wire_294, {fourFunc_wire_62_2, fourFunc_wire_103_2});
or_n #(2, 0, 0) OR_31 (fourFunc_wire_94, {fourFunc_wire_298, fourFunc_wire_296});
and_n #(2, 0, 0) AND_42 (fourFunc_wire_299, {fourFunc_wire_94_1, fourFunc_wire_300});
and_n #(2, 0, 0) AND_43 (fourFunc_wire_298, {fourFunc_wire_57_1, fourFunc_wire_99_1});
or_n #(2, 0, 0) OR_32 (fourFunc_wire_297, {fourFunc_wire_57_2, fourFunc_wire_99_2});
or_n #(2, 0, 0) OR_33 (fourFunc_wire_89, {fourFunc_wire_301, fourFunc_wire_299});
and_n #(2, 0, 0) AND_44 (fourFunc_wire_302, {fourFunc_wire_89_1, fourFunc_wire_303});
and_n #(2, 0, 0) AND_45 (fourFunc_wire_301, {fourFunc_wire_54_1, fourFunc_wire_95_1});
or_n #(2, 0, 0) OR_34 (fourFunc_wire_300, {fourFunc_wire_54_2, fourFunc_wire_95_2});
bufg #(0, 0) BUF_3 (fourFunc_wire_120, fourFunc_wire_304);
or_n #(2, 0, 0) OR_35 (fourFunc_wire_304, {fourFunc_wire_305, fourFunc_wire_302});
and_n #(2, 0, 0) AND_46 (fourFunc_wire_305, {fourFunc_wire_91_1, fourFunc_wire_90_1});
or_n #(2, 0, 0) OR_36 (fourFunc_wire_303, {fourFunc_wire_91_2, fourFunc_wire_90_2});
and_n #(2, 0, 0) AND_47 (fourFunc_wire_143, {fourFunc_wire_112, fourFunc_wire_306});
and_n #(2, 0, 0) AND_48 (fourFunc_wire_307, {fourFunc_wire_143_1, fourFunc_wire_308});
or_n #(2, 0, 0) OR_37 (fourFunc_wire_139, {fourFunc_wire_309, fourFunc_wire_307});
and_n #(2, 0, 0) AND_49 (fourFunc_wire_310, {fourFunc_wire_139_1, fourFunc_wire_311});
and_n #(2, 0, 0) AND_50 (fourFunc_wire_309, {fourFunc_wire_108_1, fourFunc_wire_144_1});
or_n #(2, 0, 0) OR_38 (fourFunc_wire_308, {fourFunc_wire_108_2, fourFunc_wire_144_2});
or_n #(2, 0, 0) OR_39 (fourFunc_wire_135, {fourFunc_wire_312, fourFunc_wire_310});
and_n #(2, 0, 0) AND_51 (fourFunc_wire_313, {fourFunc_wire_135_1, fourFunc_wire_314});
and_n #(2, 0, 0) AND_52 (fourFunc_wire_312, {fourFunc_wire_104_1, fourFunc_wire_140_1});
or_n #(2, 0, 0) OR_40 (fourFunc_wire_311, {fourFunc_wire_104_2, fourFunc_wire_140_2});
or_n #(2, 0, 0) OR_41 (fourFunc_wire_131, {fourFunc_wire_315, fourFunc_wire_313});
and_n #(2, 0, 0) AND_53 (fourFunc_wire_316, {fourFunc_wire_131_1, fourFunc_wire_317});
and_n #(2, 0, 0) AND_54 (fourFunc_wire_315, {fourFunc_wire_100_1, fourFunc_wire_136_1});
or_n #(2, 0, 0) OR_42 (fourFunc_wire_314, {fourFunc_wire_100_2, fourFunc_wire_136_2});
or_n #(2, 0, 0) OR_43 (fourFunc_wire_127, {fourFunc_wire_318, fourFunc_wire_316});
and_n #(2, 0, 0) AND_55 (fourFunc_wire_319, {fourFunc_wire_127_1, fourFunc_wire_320});
and_n #(2, 0, 0) AND_56 (fourFunc_wire_318, {fourFunc_wire_96_1, fourFunc_wire_132_1});
or_n #(2, 0, 0) OR_44 (fourFunc_wire_317, {fourFunc_wire_96_2, fourFunc_wire_132_2});
or_n #(2, 0, 0) OR_45 (fourFunc_wire_123, {fourFunc_wire_321, fourFunc_wire_319});
and_n #(2, 0, 0) AND_57 (fourFunc_wire_322, {fourFunc_wire_123_1, fourFunc_wire_323});
and_n #(2, 0, 0) AND_58 (fourFunc_wire_321, {fourFunc_wire_92_1, fourFunc_wire_128_1});
or_n #(2, 0, 0) OR_46 (fourFunc_wire_320, {fourFunc_wire_92_2, fourFunc_wire_128_2});
or_n #(2, 0, 0) OR_47 (fourFunc_wire_118, {fourFunc_wire_324, fourFunc_wire_322});
and_n #(2, 0, 0) AND_59 (fourFunc_wire_325, {fourFunc_wire_118_1, fourFunc_wire_326});
and_n #(2, 0, 0) AND_60 (fourFunc_wire_324, {fourFunc_wire_87_1, fourFunc_wire_124_1});
or_n #(2, 0, 0) OR_48 (fourFunc_wire_323, {fourFunc_wire_87_2, fourFunc_wire_124_2});
bufg #(0, 0) BUF_4 (fourFunc_wire_149, fourFunc_wire_327);
or_n #(2, 0, 0) OR_49 (fourFunc_wire_327, {fourFunc_wire_328, fourFunc_wire_325});
and_n #(2, 0, 0) AND_61 (fourFunc_wire_328, {fourFunc_wire_120_1, fourFunc_wire_119_1});
or_n #(2, 0, 0) OR_50 (fourFunc_wire_326, {fourFunc_wire_120_2, fourFunc_wire_119_2});
and_n #(2, 0, 0) AND_62 (fourFunc_wire_172, {fourFunc_wire_141, fourFunc_wire_329});
and_n #(2, 0, 0) AND_63 (fourFunc_wire_330, {fourFunc_wire_172_1, fourFunc_wire_331});
or_n #(2, 0, 0) OR_51 (fourFunc_wire_168, {fourFunc_wire_332, fourFunc_wire_330});
and_n #(2, 0, 0) AND_64 (fourFunc_wire_333, {fourFunc_wire_168_1, fourFunc_wire_334});
and_n #(2, 0, 0) AND_65 (fourFunc_wire_332, {fourFunc_wire_137_1, fourFunc_wire_173_1});
or_n #(2, 0, 0) OR_52 (fourFunc_wire_331, {fourFunc_wire_137_2, fourFunc_wire_173_2});
or_n #(2, 0, 0) OR_53 (fourFunc_wire_164, {fourFunc_wire_335, fourFunc_wire_333});
and_n #(2, 0, 0) AND_66 (fourFunc_wire_336, {fourFunc_wire_164_1, fourFunc_wire_337});
and_n #(2, 0, 0) AND_67 (fourFunc_wire_335, {fourFunc_wire_133_1, fourFunc_wire_169_1});
or_n #(2, 0, 0) OR_54 (fourFunc_wire_334, {fourFunc_wire_133_2, fourFunc_wire_169_2});
or_n #(2, 0, 0) OR_55 (fourFunc_wire_160, {fourFunc_wire_338, fourFunc_wire_336});
and_n #(2, 0, 0) AND_68 (fourFunc_wire_339, {fourFunc_wire_160_1, fourFunc_wire_340});
and_n #(2, 0, 0) AND_69 (fourFunc_wire_338, {fourFunc_wire_129_1, fourFunc_wire_165_1});
or_n #(2, 0, 0) OR_56 (fourFunc_wire_337, {fourFunc_wire_129_2, fourFunc_wire_165_2});
or_n #(2, 0, 0) OR_57 (fourFunc_wire_156, {fourFunc_wire_341, fourFunc_wire_339});
and_n #(2, 0, 0) AND_70 (fourFunc_wire_342, {fourFunc_wire_156_1, fourFunc_wire_343});
and_n #(2, 0, 0) AND_71 (fourFunc_wire_341, {fourFunc_wire_125_1, fourFunc_wire_161_1});
or_n #(2, 0, 0) OR_58 (fourFunc_wire_340, {fourFunc_wire_125_2, fourFunc_wire_161_2});
or_n #(2, 0, 0) OR_59 (fourFunc_wire_152, {fourFunc_wire_344, fourFunc_wire_342});
and_n #(2, 0, 0) AND_72 (fourFunc_wire_345, {fourFunc_wire_152_1, fourFunc_wire_346});
and_n #(2, 0, 0) AND_73 (fourFunc_wire_344, {fourFunc_wire_121_1, fourFunc_wire_157_1});
or_n #(2, 0, 0) OR_60 (fourFunc_wire_343, {fourFunc_wire_121_2, fourFunc_wire_157_2});
or_n #(2, 0, 0) OR_61 (fourFunc_wire_147, {fourFunc_wire_347, fourFunc_wire_345});
and_n #(2, 0, 0) AND_74 (fourFunc_wire_348, {fourFunc_wire_147_1, fourFunc_wire_349});
and_n #(2, 0, 0) AND_75 (fourFunc_wire_347, {fourFunc_wire_116_1, fourFunc_wire_153_1});
or_n #(2, 0, 0) OR_62 (fourFunc_wire_346, {fourFunc_wire_116_2, fourFunc_wire_153_2});
bufg #(0, 0) BUF_5 (fourFunc_wire_178, fourFunc_wire_350);
or_n #(2, 0, 0) OR_63 (fourFunc_wire_350, {fourFunc_wire_351, fourFunc_wire_348});
and_n #(2, 0, 0) AND_76 (fourFunc_wire_351, {fourFunc_wire_149_1, fourFunc_wire_148_1});
or_n #(2, 0, 0) OR_64 (fourFunc_wire_349, {fourFunc_wire_149_2, fourFunc_wire_148_2});
and_n #(2, 0, 0) AND_77 (fourFunc_wire_201, {fourFunc_wire_170, fourFunc_wire_352});
and_n #(2, 0, 0) AND_78 (fourFunc_wire_353, {fourFunc_wire_201_1, fourFunc_wire_354});
or_n #(2, 0, 0) OR_65 (fourFunc_wire_197, {fourFunc_wire_355, fourFunc_wire_353});
and_n #(2, 0, 0) AND_79 (fourFunc_wire_356, {fourFunc_wire_197_1, fourFunc_wire_357});
and_n #(2, 0, 0) AND_80 (fourFunc_wire_355, {fourFunc_wire_166_1, fourFunc_wire_202_1});
or_n #(2, 0, 0) OR_66 (fourFunc_wire_354, {fourFunc_wire_166_2, fourFunc_wire_202_2});
or_n #(2, 0, 0) OR_67 (fourFunc_wire_193, {fourFunc_wire_358, fourFunc_wire_356});
and_n #(2, 0, 0) AND_81 (fourFunc_wire_359, {fourFunc_wire_193_1, fourFunc_wire_360});
and_n #(2, 0, 0) AND_82 (fourFunc_wire_358, {fourFunc_wire_162_1, fourFunc_wire_198_1});
or_n #(2, 0, 0) OR_68 (fourFunc_wire_357, {fourFunc_wire_162_2, fourFunc_wire_198_2});
or_n #(2, 0, 0) OR_69 (fourFunc_wire_189, {fourFunc_wire_361, fourFunc_wire_359});
and_n #(2, 0, 0) AND_83 (fourFunc_wire_362, {fourFunc_wire_189_1, fourFunc_wire_363});
and_n #(2, 0, 0) AND_84 (fourFunc_wire_361, {fourFunc_wire_158_1, fourFunc_wire_194_1});
or_n #(2, 0, 0) OR_70 (fourFunc_wire_360, {fourFunc_wire_158_2, fourFunc_wire_194_2});
or_n #(2, 0, 0) OR_71 (fourFunc_wire_185, {fourFunc_wire_364, fourFunc_wire_362});
and_n #(2, 0, 0) AND_85 (fourFunc_wire_365, {fourFunc_wire_185_1, fourFunc_wire_366});
and_n #(2, 0, 0) AND_86 (fourFunc_wire_364, {fourFunc_wire_154_1, fourFunc_wire_190_1});
or_n #(2, 0, 0) OR_72 (fourFunc_wire_363, {fourFunc_wire_154_2, fourFunc_wire_190_2});
or_n #(2, 0, 0) OR_73 (fourFunc_wire_181, {fourFunc_wire_367, fourFunc_wire_365});
and_n #(2, 0, 0) AND_87 (fourFunc_wire_368, {fourFunc_wire_181_1, fourFunc_wire_369});
and_n #(2, 0, 0) AND_88 (fourFunc_wire_367, {fourFunc_wire_150_1, fourFunc_wire_186_1});
or_n #(2, 0, 0) OR_74 (fourFunc_wire_366, {fourFunc_wire_150_2, fourFunc_wire_186_2});
or_n #(2, 0, 0) OR_75 (fourFunc_wire_176, {fourFunc_wire_370, fourFunc_wire_368});
and_n #(2, 0, 0) AND_89 (fourFunc_wire_371, {fourFunc_wire_176_1, fourFunc_wire_372});
and_n #(2, 0, 0) AND_90 (fourFunc_wire_370, {fourFunc_wire_145_1, fourFunc_wire_182_1});
or_n #(2, 0, 0) OR_76 (fourFunc_wire_369, {fourFunc_wire_145_2, fourFunc_wire_182_2});
bufg #(0, 0) BUF_6 (fourFunc_wire_207, fourFunc_wire_373);
or_n #(2, 0, 0) OR_77 (fourFunc_wire_373, {fourFunc_wire_374, fourFunc_wire_371});
and_n #(2, 0, 0) AND_91 (fourFunc_wire_374, {fourFunc_wire_178_1, fourFunc_wire_177_1});
or_n #(2, 0, 0) OR_78 (fourFunc_wire_372, {fourFunc_wire_178_2, fourFunc_wire_177_2});
and_n #(2, 0, 0) AND_92 (fourFunc_wire_230, {fourFunc_wire_199, fourFunc_wire_375});
and_n #(2, 0, 0) AND_93 (fourFunc_wire_376, {fourFunc_wire_230_1, fourFunc_wire_377});
or_n #(2, 0, 0) OR_79 (fourFunc_wire_226, {fourFunc_wire_378, fourFunc_wire_376});
and_n #(2, 0, 0) AND_94 (fourFunc_wire_379, {fourFunc_wire_226_1, fourFunc_wire_380});
and_n #(2, 0, 0) AND_95 (fourFunc_wire_378, {fourFunc_wire_195_1, fourFunc_wire_231_1});
or_n #(2, 0, 0) OR_80 (fourFunc_wire_377, {fourFunc_wire_195_2, fourFunc_wire_231_2});
or_n #(2, 0, 0) OR_81 (fourFunc_wire_222, {fourFunc_wire_381, fourFunc_wire_379});
and_n #(2, 0, 0) AND_96 (fourFunc_wire_382, {fourFunc_wire_222_1, fourFunc_wire_383});
and_n #(2, 0, 0) AND_97 (fourFunc_wire_381, {fourFunc_wire_191_1, fourFunc_wire_227_1});
or_n #(2, 0, 0) OR_82 (fourFunc_wire_380, {fourFunc_wire_191_2, fourFunc_wire_227_2});
or_n #(2, 0, 0) OR_83 (fourFunc_wire_218, {fourFunc_wire_384, fourFunc_wire_382});
and_n #(2, 0, 0) AND_98 (fourFunc_wire_385, {fourFunc_wire_218_1, fourFunc_wire_386});
and_n #(2, 0, 0) AND_99 (fourFunc_wire_384, {fourFunc_wire_187_1, fourFunc_wire_223_1});
or_n #(2, 0, 0) OR_84 (fourFunc_wire_383, {fourFunc_wire_187_2, fourFunc_wire_223_2});
or_n #(2, 0, 0) OR_85 (fourFunc_wire_214, {fourFunc_wire_387, fourFunc_wire_385});
and_n #(2, 0, 0) AND_100 (fourFunc_wire_388, {fourFunc_wire_214_1, fourFunc_wire_389});
and_n #(2, 0, 0) AND_101 (fourFunc_wire_387, {fourFunc_wire_183_1, fourFunc_wire_219_1});
or_n #(2, 0, 0) OR_86 (fourFunc_wire_386, {fourFunc_wire_183_2, fourFunc_wire_219_2});
or_n #(2, 0, 0) OR_87 (fourFunc_wire_210, {fourFunc_wire_390, fourFunc_wire_388});
and_n #(2, 0, 0) AND_102 (fourFunc_wire_391, {fourFunc_wire_210_1, fourFunc_wire_392});
and_n #(2, 0, 0) AND_103 (fourFunc_wire_390, {fourFunc_wire_179_1, fourFunc_wire_215_1});
or_n #(2, 0, 0) OR_88 (fourFunc_wire_389, {fourFunc_wire_179_2, fourFunc_wire_215_2});
or_n #(2, 0, 0) OR_89 (fourFunc_wire_205, {fourFunc_wire_393, fourFunc_wire_391});
and_n #(2, 0, 0) AND_104 (fourFunc_wire_394, {fourFunc_wire_205_1, fourFunc_wire_395});
and_n #(2, 0, 0) AND_105 (fourFunc_wire_393, {fourFunc_wire_174_1, fourFunc_wire_211_1});
or_n #(2, 0, 0) OR_90 (fourFunc_wire_392, {fourFunc_wire_174_2, fourFunc_wire_211_2});
bufg #(0, 0) BUF_7 (fourFunc_wire_236, fourFunc_wire_396);
or_n #(2, 0, 0) OR_91 (fourFunc_wire_396, {fourFunc_wire_397, fourFunc_wire_394});
and_n #(2, 0, 0) AND_106 (fourFunc_wire_397, {fourFunc_wire_207_1, fourFunc_wire_206_1});
or_n #(2, 0, 0) OR_92 (fourFunc_wire_395, {fourFunc_wire_207_2, fourFunc_wire_206_2});
and_n #(2, 0, 0) AND_107 (fourFunc_wire_259, {fourFunc_wire_228, fourFunc_wire_398});
and_n #(2, 0, 0) AND_108 (fourFunc_wire_399, {fourFunc_wire_259_1, fourFunc_wire_400});
or_n #(2, 0, 0) OR_93 (fourFunc_wire_255, {fourFunc_wire_401, fourFunc_wire_399});
and_n #(2, 0, 0) AND_109 (fourFunc_wire_402, {fourFunc_wire_255_1, fourFunc_wire_403});
and_n #(2, 0, 0) AND_110 (fourFunc_wire_401, {fourFunc_wire_224_1, fourFunc_wire_260_1});
or_n #(2, 0, 0) OR_94 (fourFunc_wire_400, {fourFunc_wire_224_2, fourFunc_wire_260_2});
or_n #(2, 0, 0) OR_95 (fourFunc_wire_251, {fourFunc_wire_404, fourFunc_wire_402});
and_n #(2, 0, 0) AND_111 (fourFunc_wire_405, {fourFunc_wire_251_1, fourFunc_wire_406});
and_n #(2, 0, 0) AND_112 (fourFunc_wire_404, {fourFunc_wire_220_1, fourFunc_wire_256_1});
or_n #(2, 0, 0) OR_96 (fourFunc_wire_403, {fourFunc_wire_220_2, fourFunc_wire_256_2});
or_n #(2, 0, 0) OR_97 (fourFunc_wire_247, {fourFunc_wire_407, fourFunc_wire_405});
and_n #(2, 0, 0) AND_113 (fourFunc_wire_408, {fourFunc_wire_247_1, fourFunc_wire_409});
and_n #(2, 0, 0) AND_114 (fourFunc_wire_407, {fourFunc_wire_216_1, fourFunc_wire_252_1});
or_n #(2, 0, 0) OR_98 (fourFunc_wire_406, {fourFunc_wire_216_2, fourFunc_wire_252_2});
or_n #(2, 0, 0) OR_99 (fourFunc_wire_243, {fourFunc_wire_410, fourFunc_wire_408});
and_n #(2, 0, 0) AND_115 (fourFunc_wire_411, {fourFunc_wire_243_1, fourFunc_wire_412});
and_n #(2, 0, 0) AND_116 (fourFunc_wire_410, {fourFunc_wire_212_1, fourFunc_wire_248_1});
or_n #(2, 0, 0) OR_100 (fourFunc_wire_409, {fourFunc_wire_212_2, fourFunc_wire_248_2});
or_n #(2, 0, 0) OR_101 (fourFunc_wire_239, {fourFunc_wire_413, fourFunc_wire_411});
and_n #(2, 0, 0) AND_117 (fourFunc_wire_414, {fourFunc_wire_239_1, fourFunc_wire_415});
and_n #(2, 0, 0) AND_118 (fourFunc_wire_413, {fourFunc_wire_208_1, fourFunc_wire_244_1});
or_n #(2, 0, 0) OR_102 (fourFunc_wire_412, {fourFunc_wire_208_2, fourFunc_wire_244_2});
or_n #(2, 0, 0) OR_103 (fourFunc_wire_234, {fourFunc_wire_416, fourFunc_wire_414});
and_n #(2, 0, 0) AND_119 (fourFunc_wire_417, {fourFunc_wire_234_1, fourFunc_wire_418});
and_n #(2, 0, 0) AND_120 (fourFunc_wire_416, {fourFunc_wire_203_1, fourFunc_wire_240_1});
or_n #(2, 0, 0) OR_104 (fourFunc_wire_415, {fourFunc_wire_203_2, fourFunc_wire_240_2});
bufg #(0, 0) BUF_8 (fourFunc_wire_419, fourFunc_wire_420);
or_n #(2, 0, 0) OR_105 (fourFunc_wire_420, {fourFunc_wire_421, fourFunc_wire_417});
and_n #(2, 0, 0) AND_121 (fourFunc_wire_421, {fourFunc_wire_236_1, fourFunc_wire_235_1});
or_n #(2, 0, 0) OR_106 (fourFunc_wire_418, {fourFunc_wire_236_2, fourFunc_wire_235_2});
and_n #(2, 0, 0) AND_122 (fourFunc_wire_61, {fourFunc_wire_422_0, fourFunc_wire_423_0});
and_n #(2, 0, 0) AND_123 (fourFunc_wire_66, {fourFunc_wire_422_1, fourFunc_wire_424_0});
and_n #(2, 0, 0) AND_124 (fourFunc_wire_71, {fourFunc_wire_422_2, fourFunc_wire_425_0});
and_n #(2, 0, 0) AND_125 (fourFunc_wire_76, {fourFunc_wire_422_3, fourFunc_wire_426_0});
and_n #(2, 0, 0) AND_126 (fourFunc_wire_81, {fourFunc_wire_422_4, fourFunc_wire_427_0});
and_n #(2, 0, 0) AND_127 (fourFunc_wire_86, {fourFunc_wire_422_5, fourFunc_wire_428_0});
and_n #(2, 0, 0) AND_128 (fourFunc_wire_262, {fourFunc_wire_422_6, fourFunc_wire_429_0});
and_n #(2, 0, 0) AND_129 (fourFunc_wire_261, {fourFunc_wire_430_0, fourFunc_wire_423_1});
and_n #(2, 0, 0) AND_130 (fourFunc_wire_60, {fourFunc_wire_430_1, fourFunc_wire_424_1});
and_n #(2, 0, 0) AND_131 (fourFunc_wire_65, {fourFunc_wire_430_2, fourFunc_wire_425_1});
and_n #(2, 0, 0) AND_132 (fourFunc_wire_70, {fourFunc_wire_430_3, fourFunc_wire_426_1});
and_n #(2, 0, 0) AND_133 (fourFunc_wire_75, {fourFunc_wire_430_4, fourFunc_wire_427_1});
and_n #(2, 0, 0) AND_134 (fourFunc_wire_80, {fourFunc_wire_430_5, fourFunc_wire_428_1});
and_n #(2, 0, 0) AND_135 (fourFunc_wire_85, {fourFunc_wire_430_6, fourFunc_wire_429_1});
and_n #(2, 0, 0) AND_136 (fourFunc_wire_263, {fourFunc_wire_430_7, fourFunc_wire_431_0});
and_n #(2, 0, 0) AND_137 (fourFunc_wire_90, {fourFunc_wire_432_0, fourFunc_wire_423_2});
and_n #(2, 0, 0) AND_138 (fourFunc_wire_95, {fourFunc_wire_432_1, fourFunc_wire_424_2});
and_n #(2, 0, 0) AND_139 (fourFunc_wire_99, {fourFunc_wire_432_2, fourFunc_wire_425_2});
and_n #(2, 0, 0) AND_140 (fourFunc_wire_103, {fourFunc_wire_432_3, fourFunc_wire_426_2});
and_n #(2, 0, 0) AND_141 (fourFunc_wire_107, {fourFunc_wire_432_4, fourFunc_wire_427_2});
and_n #(2, 0, 0) AND_142 (fourFunc_wire_111, {fourFunc_wire_432_5, fourFunc_wire_428_2});
and_n #(2, 0, 0) AND_143 (fourFunc_wire_115, {fourFunc_wire_432_6, fourFunc_wire_429_2});
and_n #(2, 0, 0) AND_144 (fourFunc_wire_283, {fourFunc_wire_432_7, fourFunc_wire_431_1});
and_n #(2, 0, 0) AND_145 (fourFunc_wire_119, {fourFunc_wire_433_0, fourFunc_wire_423_3});
and_n #(2, 0, 0) AND_146 (fourFunc_wire_124, {fourFunc_wire_433_1, fourFunc_wire_424_3});
and_n #(2, 0, 0) AND_147 (fourFunc_wire_128, {fourFunc_wire_433_2, fourFunc_wire_425_3});
and_n #(2, 0, 0) AND_148 (fourFunc_wire_132, {fourFunc_wire_433_3, fourFunc_wire_426_3});
and_n #(2, 0, 0) AND_149 (fourFunc_wire_136, {fourFunc_wire_433_4, fourFunc_wire_427_3});
and_n #(2, 0, 0) AND_150 (fourFunc_wire_140, {fourFunc_wire_433_5, fourFunc_wire_428_3});
and_n #(2, 0, 0) AND_151 (fourFunc_wire_144, {fourFunc_wire_433_6, fourFunc_wire_429_3});
and_n #(2, 0, 0) AND_152 (fourFunc_wire_306, {fourFunc_wire_433_7, fourFunc_wire_431_2});
and_n #(2, 0, 0) AND_153 (fourFunc_wire_148, {fourFunc_wire_434_0, fourFunc_wire_423_4});
and_n #(2, 0, 0) AND_154 (fourFunc_wire_153, {fourFunc_wire_434_1, fourFunc_wire_424_4});
and_n #(2, 0, 0) AND_155 (fourFunc_wire_157, {fourFunc_wire_434_2, fourFunc_wire_425_4});
and_n #(2, 0, 0) AND_156 (fourFunc_wire_161, {fourFunc_wire_434_3, fourFunc_wire_426_4});
and_n #(2, 0, 0) AND_157 (fourFunc_wire_165, {fourFunc_wire_434_4, fourFunc_wire_427_4});
and_n #(2, 0, 0) AND_158 (fourFunc_wire_169, {fourFunc_wire_434_5, fourFunc_wire_428_4});
and_n #(2, 0, 0) AND_159 (fourFunc_wire_173, {fourFunc_wire_434_6, fourFunc_wire_429_4});
and_n #(2, 0, 0) AND_160 (fourFunc_wire_329, {fourFunc_wire_434_7, fourFunc_wire_431_3});
and_n #(2, 0, 0) AND_161 (fourFunc_wire_177, {fourFunc_wire_435_0, fourFunc_wire_423_5});
and_n #(2, 0, 0) AND_162 (fourFunc_wire_182, {fourFunc_wire_435_1, fourFunc_wire_424_5});
and_n #(2, 0, 0) AND_163 (fourFunc_wire_186, {fourFunc_wire_435_2, fourFunc_wire_425_5});
and_n #(2, 0, 0) AND_164 (fourFunc_wire_190, {fourFunc_wire_435_3, fourFunc_wire_426_5});
and_n #(2, 0, 0) AND_165 (fourFunc_wire_194, {fourFunc_wire_435_4, fourFunc_wire_427_5});
and_n #(2, 0, 0) AND_166 (fourFunc_wire_198, {fourFunc_wire_435_5, fourFunc_wire_428_5});
and_n #(2, 0, 0) AND_167 (fourFunc_wire_202, {fourFunc_wire_435_6, fourFunc_wire_429_5});
and_n #(2, 0, 0) AND_168 (fourFunc_wire_352, {fourFunc_wire_435_7, fourFunc_wire_431_4});
and_n #(2, 0, 0) AND_169 (fourFunc_wire_206, {fourFunc_wire_436_0, fourFunc_wire_423_6});
and_n #(2, 0, 0) AND_170 (fourFunc_wire_211, {fourFunc_wire_436_1, fourFunc_wire_424_6});
and_n #(2, 0, 0) AND_171 (fourFunc_wire_215, {fourFunc_wire_436_2, fourFunc_wire_425_6});
and_n #(2, 0, 0) AND_172 (fourFunc_wire_219, {fourFunc_wire_436_3, fourFunc_wire_426_6});
and_n #(2, 0, 0) AND_173 (fourFunc_wire_223, {fourFunc_wire_436_4, fourFunc_wire_427_6});
and_n #(2, 0, 0) AND_174 (fourFunc_wire_227, {fourFunc_wire_436_5, fourFunc_wire_428_6});
and_n #(2, 0, 0) AND_175 (fourFunc_wire_231, {fourFunc_wire_436_6, fourFunc_wire_429_6});
and_n #(2, 0, 0) AND_176 (fourFunc_wire_375, {fourFunc_wire_436_7, fourFunc_wire_431_5});
and_n #(2, 0, 0) AND_177 (fourFunc_wire_235, {fourFunc_wire_437_0, fourFunc_wire_423_7});
and_n #(2, 0, 0) AND_178 (fourFunc_wire_240, {fourFunc_wire_437_1, fourFunc_wire_424_7});
and_n #(2, 0, 0) AND_179 (fourFunc_wire_244, {fourFunc_wire_437_2, fourFunc_wire_425_7});
and_n #(2, 0, 0) AND_180 (fourFunc_wire_248, {fourFunc_wire_437_3, fourFunc_wire_426_7});
and_n #(2, 0, 0) AND_181 (fourFunc_wire_252, {fourFunc_wire_437_4, fourFunc_wire_427_7});
and_n #(2, 0, 0) AND_182 (fourFunc_wire_256, {fourFunc_wire_437_5, fourFunc_wire_428_7});
and_n #(2, 0, 0) AND_183 (fourFunc_wire_260, {fourFunc_wire_437_6, fourFunc_wire_429_7});
and_n #(2, 0, 0) AND_184 (fourFunc_wire_398, {fourFunc_wire_437_7, fourFunc_wire_431_6});
xor_n #(2, 0, 0) XOR_98 (fourFunc_wire_438, {fourFunc_wire_439, fourFunc_wire_3_11});
xor_n #(2, 0, 0) XOR_99 (fourFunc_wire_440, {fourFunc_wire_11_9, fourFunc_wire_2_15});
xnor_n #(2, 0, 0) XNOR_1 (fourFunc_wire_441, {fourFunc_wire_422_7, fourFunc_wire_442_0});
xnor_n #(2, 0, 0) XNOR_2 (fourFunc_wire_443, {fourFunc_wire_444_0, fourFunc_wire_445});
xnor_n #(2, 0, 0) XNOR_3 (fourFunc_wire_446, {fourFunc_wire_447_0, fourFunc_wire_448_0});
xor_n #(2, 0, 0) XOR_100 (fourFunc_wire_449, {fourFunc_wire_450, fourFunc_wire_451_0});
xnor_n #(2, 0, 0) XNOR_4 (fourFunc_wire_450, {fourFunc_wire_452_0, fourFunc_wire_437_8});
xor_n #(2, 0, 0) XOR_101 (fourFunc_wire_453, {fourFunc_wire_454, fourFunc_wire_455_0});
xnor_n #(2, 0, 0) XNOR_5 (fourFunc_wire_454, {fourFunc_wire_456_0, fourFunc_wire_436_8});
xor_n #(2, 0, 0) XOR_102 (fourFunc_wire_457, {fourFunc_wire_458, fourFunc_wire_459_0});
xnor_n #(2, 0, 0) XNOR_6 (fourFunc_wire_458, {fourFunc_wire_460_0, fourFunc_wire_435_8});
xor_n #(2, 0, 0) XOR_103 (fourFunc_wire_461, {fourFunc_wire_462, fourFunc_wire_463_0});
xnor_n #(2, 0, 0) XNOR_7 (fourFunc_wire_462, {fourFunc_wire_464_0, fourFunc_wire_434_8});
xor_n #(2, 0, 0) XOR_104 (fourFunc_wire_465, {fourFunc_wire_466, fourFunc_wire_467_0});
xnor_n #(2, 0, 0) XNOR_8 (fourFunc_wire_466, {fourFunc_wire_468_0, fourFunc_wire_433_8});
xor_n #(2, 0, 0) XOR_105 (fourFunc_wire_469, {fourFunc_wire_470, fourFunc_wire_471_0});
xnor_n #(2, 0, 0) XNOR_9 (fourFunc_wire_470, {fourFunc_wire_472_0, fourFunc_wire_432_8});
xor_n #(2, 0, 0) XOR_106 (fourFunc_wire_473, {fourFunc_wire_474, fourFunc_wire_475_0});
xnor_n #(2, 0, 0) XNOR_10 (fourFunc_wire_474, {fourFunc_wire_476_0, fourFunc_wire_430_8});
xor_n #(2, 0, 0) XOR_107 (fourFunc_wire_477, {fourFunc_wire_442_1, fourFunc_wire_422_8});
xor_n #(2, 0, 0) XOR_108 (fourFunc_wire_478, {fourFunc_wire_479_0, fourFunc_wire_447_1});
xor_n #(2, 0, 0) XOR_109 (fourFunc_wire_480, {fourFunc_wire_481, fourFunc_wire_444_1});
xor_n #(2, 0, 0) XOR_110 (fourFunc_wire_482, {fourFunc_wire_483, fourFunc_wire_484_0});
xor_n #(2, 0, 0) XOR_111 (fourFunc_wire_483, {fourFunc_wire_437_9, fourFunc_wire_452_1});
xor_n #(2, 0, 0) XOR_112 (fourFunc_wire_485, {fourFunc_wire_486, fourFunc_wire_487_0});
xor_n #(2, 0, 0) XOR_113 (fourFunc_wire_486, {fourFunc_wire_436_9, fourFunc_wire_456_1});
xor_n #(2, 0, 0) XOR_114 (fourFunc_wire_488, {fourFunc_wire_489, fourFunc_wire_490_0});
xor_n #(2, 0, 0) XOR_115 (fourFunc_wire_489, {fourFunc_wire_435_9, fourFunc_wire_460_1});
xor_n #(2, 0, 0) XOR_116 (fourFunc_wire_491, {fourFunc_wire_492, fourFunc_wire_493_0});
xor_n #(2, 0, 0) XOR_117 (fourFunc_wire_492, {fourFunc_wire_434_9, fourFunc_wire_464_1});
xor_n #(2, 0, 0) XOR_118 (fourFunc_wire_494, {fourFunc_wire_495, fourFunc_wire_496_0});
xor_n #(2, 0, 0) XOR_119 (fourFunc_wire_495, {fourFunc_wire_433_9, fourFunc_wire_468_1});
xor_n #(2, 0, 0) XOR_120 (fourFunc_wire_497, {fourFunc_wire_498, fourFunc_wire_499_0});
xor_n #(2, 0, 0) XOR_121 (fourFunc_wire_498, {fourFunc_wire_432_9, fourFunc_wire_472_1});
xor_n #(2, 0, 0) XOR_122 (fourFunc_wire_500, {fourFunc_wire_501, fourFunc_wire_502_0});
xor_n #(2, 0, 0) XOR_123 (fourFunc_wire_501, {fourFunc_wire_430_9, fourFunc_wire_476_1});
and_n #(2, 0, 0) AND_185 (fourFunc_wire_502, {fourFunc_wire_442_2, fourFunc_wire_422_9});
and_n #(2, 0, 0) AND_186 (fourFunc_wire_503, {fourFunc_wire_502_1, fourFunc_wire_504});
and_n #(2, 0, 0) AND_187 (fourFunc_wire_481, {fourFunc_wire_479_1, fourFunc_wire_447_2});
or_n #(2, 0, 0) OR_107 (fourFunc_wire_499, {fourFunc_wire_505, fourFunc_wire_503});
and_n #(2, 0, 0) AND_188 (fourFunc_wire_506, {fourFunc_wire_499_1, fourFunc_wire_507});
and_n #(2, 0, 0) AND_189 (fourFunc_wire_505, {fourFunc_wire_476_2, fourFunc_wire_430_10});
or_n #(2, 0, 0) OR_108 (fourFunc_wire_504, {fourFunc_wire_476_3, fourFunc_wire_430_11});
or_n #(2, 0, 0) OR_109 (fourFunc_wire_496, {fourFunc_wire_508, fourFunc_wire_506});
and_n #(2, 0, 0) AND_190 (fourFunc_wire_509, {fourFunc_wire_496_1, fourFunc_wire_510});
and_n #(2, 0, 0) AND_191 (fourFunc_wire_508, {fourFunc_wire_472_2, fourFunc_wire_432_10});
or_n #(2, 0, 0) OR_110 (fourFunc_wire_507, {fourFunc_wire_472_3, fourFunc_wire_432_11});
or_n #(2, 0, 0) OR_111 (fourFunc_wire_493, {fourFunc_wire_511, fourFunc_wire_509});
and_n #(2, 0, 0) AND_192 (fourFunc_wire_512, {fourFunc_wire_493_1, fourFunc_wire_513});
and_n #(2, 0, 0) AND_193 (fourFunc_wire_511, {fourFunc_wire_468_2, fourFunc_wire_433_10});
or_n #(2, 0, 0) OR_112 (fourFunc_wire_510, {fourFunc_wire_468_3, fourFunc_wire_433_11});
or_n #(2, 0, 0) OR_113 (fourFunc_wire_490, {fourFunc_wire_514, fourFunc_wire_512});
and_n #(2, 0, 0) AND_194 (fourFunc_wire_515, {fourFunc_wire_490_1, fourFunc_wire_516});
and_n #(2, 0, 0) AND_195 (fourFunc_wire_514, {fourFunc_wire_464_2, fourFunc_wire_434_10});
or_n #(2, 0, 0) OR_114 (fourFunc_wire_513, {fourFunc_wire_464_3, fourFunc_wire_434_11});
or_n #(2, 0, 0) OR_115 (fourFunc_wire_487, {fourFunc_wire_517, fourFunc_wire_515});
and_n #(2, 0, 0) AND_196 (fourFunc_wire_518, {fourFunc_wire_487_1, fourFunc_wire_519});
and_n #(2, 0, 0) AND_197 (fourFunc_wire_517, {fourFunc_wire_460_2, fourFunc_wire_435_10});
or_n #(2, 0, 0) OR_116 (fourFunc_wire_516, {fourFunc_wire_460_3, fourFunc_wire_435_11});
or_n #(2, 0, 0) OR_117 (fourFunc_wire_484, {fourFunc_wire_520, fourFunc_wire_518});
and_n #(2, 0, 0) AND_198 (fourFunc_wire_521, {fourFunc_wire_484_1, fourFunc_wire_522});
and_n #(2, 0, 0) AND_199 (fourFunc_wire_520, {fourFunc_wire_456_2, fourFunc_wire_436_10});
or_n #(2, 0, 0) OR_118 (fourFunc_wire_519, {fourFunc_wire_456_3, fourFunc_wire_436_11});
or_n #(2, 0, 0) OR_119 (fourFunc_wire_479, {fourFunc_wire_523, fourFunc_wire_521});
and_n #(2, 0, 0) AND_200 (fourFunc_wire_523, {fourFunc_wire_452_2, fourFunc_wire_437_10});
or_n #(2, 0, 0) OR_120 (fourFunc_wire_522, {fourFunc_wire_452_3, fourFunc_wire_437_11});
or_n #(2, 0, 0) OR_121 (fourFunc_wire_475, {fourFunc_wire_524, fourFunc_wire_442_3});
and_n #(2, 0, 0) AND_201 (fourFunc_wire_525, {fourFunc_wire_475_1, fourFunc_wire_526});
notg #(0, 0) NOT_15 (fourFunc_wire_524, fourFunc_wire_422_10);
or_n #(2, 0, 0) OR_122 (fourFunc_wire_471, {fourFunc_wire_527, fourFunc_wire_525});
and_n #(2, 0, 0) AND_202 (fourFunc_wire_528, {fourFunc_wire_471_1, fourFunc_wire_529});
notg #(0, 0) NOT_16 (fourFunc_wire_530, fourFunc_wire_430_12);
or_n #(2, 0, 0) OR_123 (fourFunc_wire_526, {fourFunc_wire_530, fourFunc_wire_476_4});
notg #(0, 0) NOT_17 (fourFunc_wire_531, fourFunc_wire_430_13);
and_n #(2, 0, 0) AND_203 (fourFunc_wire_527, {fourFunc_wire_531, fourFunc_wire_476_5});
or_n #(2, 0, 0) OR_124 (fourFunc_wire_467, {fourFunc_wire_532, fourFunc_wire_528});
and_n #(2, 0, 0) AND_204 (fourFunc_wire_533, {fourFunc_wire_467_1, fourFunc_wire_534});
notg #(0, 0) NOT_18 (fourFunc_wire_535, fourFunc_wire_432_12);
or_n #(2, 0, 0) OR_125 (fourFunc_wire_529, {fourFunc_wire_535, fourFunc_wire_472_4});
notg #(0, 0) NOT_19 (fourFunc_wire_536, fourFunc_wire_432_13);
and_n #(2, 0, 0) AND_205 (fourFunc_wire_532, {fourFunc_wire_536, fourFunc_wire_472_5});
or_n #(2, 0, 0) OR_126 (fourFunc_wire_463, {fourFunc_wire_537, fourFunc_wire_533});
and_n #(2, 0, 0) AND_206 (fourFunc_wire_538, {fourFunc_wire_463_1, fourFunc_wire_539});
notg #(0, 0) NOT_20 (fourFunc_wire_540, fourFunc_wire_433_12);
or_n #(2, 0, 0) OR_127 (fourFunc_wire_534, {fourFunc_wire_540, fourFunc_wire_468_4});
notg #(0, 0) NOT_21 (fourFunc_wire_541, fourFunc_wire_433_13);
and_n #(2, 0, 0) AND_207 (fourFunc_wire_537, {fourFunc_wire_541, fourFunc_wire_468_5});
or_n #(2, 0, 0) OR_128 (fourFunc_wire_459, {fourFunc_wire_542, fourFunc_wire_538});
and_n #(2, 0, 0) AND_208 (fourFunc_wire_543, {fourFunc_wire_459_1, fourFunc_wire_544});
notg #(0, 0) NOT_22 (fourFunc_wire_545, fourFunc_wire_434_12);
or_n #(2, 0, 0) OR_129 (fourFunc_wire_539, {fourFunc_wire_545, fourFunc_wire_464_4});
notg #(0, 0) NOT_23 (fourFunc_wire_546, fourFunc_wire_434_13);
and_n #(2, 0, 0) AND_209 (fourFunc_wire_542, {fourFunc_wire_546, fourFunc_wire_464_5});
or_n #(2, 0, 0) OR_130 (fourFunc_wire_455, {fourFunc_wire_547, fourFunc_wire_543});
and_n #(2, 0, 0) AND_210 (fourFunc_wire_548, {fourFunc_wire_455_1, fourFunc_wire_549});
notg #(0, 0) NOT_24 (fourFunc_wire_550, fourFunc_wire_435_12);
or_n #(2, 0, 0) OR_131 (fourFunc_wire_544, {fourFunc_wire_550, fourFunc_wire_460_4});
notg #(0, 0) NOT_25 (fourFunc_wire_551, fourFunc_wire_435_13);
and_n #(2, 0, 0) AND_211 (fourFunc_wire_547, {fourFunc_wire_551, fourFunc_wire_460_5});
or_n #(2, 0, 0) OR_132 (fourFunc_wire_451, {fourFunc_wire_552, fourFunc_wire_548});
and_n #(2, 0, 0) AND_212 (fourFunc_wire_553, {fourFunc_wire_451_1, fourFunc_wire_554});
notg #(0, 0) NOT_26 (fourFunc_wire_555, fourFunc_wire_436_12);
or_n #(2, 0, 0) OR_133 (fourFunc_wire_549, {fourFunc_wire_555, fourFunc_wire_456_4});
notg #(0, 0) NOT_27 (fourFunc_wire_556, fourFunc_wire_436_13);
and_n #(2, 0, 0) AND_213 (fourFunc_wire_552, {fourFunc_wire_556, fourFunc_wire_456_5});
and_n #(2, 0, 0) AND_214 (fourFunc_wire_557, {fourFunc_wire_448_1, fourFunc_wire_447_3});
or_n #(3, 0, 0) OR_134 (fourFunc_wire_445, {fourFunc_wire_448_2, fourFunc_wire_557, fourFunc_wire_447_4});
or_n #(2, 0, 0) OR_135 (fourFunc_wire_448, {fourFunc_wire_558, fourFunc_wire_553});
notg #(0, 0) NOT_28 (fourFunc_wire_559, fourFunc_wire_437_12);
or_n #(2, 0, 0) OR_136 (fourFunc_wire_554, {fourFunc_wire_559, fourFunc_wire_452_4});
notg #(0, 0) NOT_29 (fourFunc_wire_560, fourFunc_wire_437_13);
and_n #(2, 0, 0) AND_215 (fourFunc_wire_558, {fourFunc_wire_560, fourFunc_wire_452_5});
bufg #(0, 0) BUF_9 (fourFunc_wire_561, 1'b0);
and_n #(2, 0, 0) AND_216 (fourFunc_wire_572, {fourFunc_wire_477, fourFunc_wire_563_0});
and_n #(2, 0, 0) AND_217 (fourFunc_wire_573, {fourFunc_wire_500, fourFunc_wire_563_1});
and_n #(2, 0, 0) AND_218 (fourFunc_wire_574, {fourFunc_wire_497, fourFunc_wire_563_2});
and_n #(2, 0, 0) AND_219 (fourFunc_wire_575, {fourFunc_wire_494, fourFunc_wire_563_3});
and_n #(2, 0, 0) AND_220 (fourFunc_wire_576, {fourFunc_wire_491, fourFunc_wire_563_4});
and_n #(2, 0, 0) AND_221 (fourFunc_wire_577, {fourFunc_wire_488, fourFunc_wire_563_5});
and_n #(2, 0, 0) AND_222 (fourFunc_wire_578, {fourFunc_wire_485, fourFunc_wire_563_6});
and_n #(2, 0, 0) AND_223 (fourFunc_wire_579, {fourFunc_wire_482, fourFunc_wire_563_7});
and_n #(2, 0, 0) AND_224 (fourFunc_wire_580, {fourFunc_wire_478, fourFunc_wire_563_8});
and_n #(2, 0, 0) AND_225 (fourFunc_wire_581, {fourFunc_wire_480, fourFunc_wire_563_9});
notg #(0, 0) NOT_30 (fourFunc_wire_582, fourFunc_wire_563_10);
notg #(0, 0) NOT_31 (fourFunc_wire_583, fourFunc_wire_563_11);
notg #(0, 0) NOT_32 (fourFunc_wire_584, fourFunc_wire_563_12);
notg #(0, 0) NOT_33 (fourFunc_wire_585, fourFunc_wire_563_13);
notg #(0, 0) NOT_34 (fourFunc_wire_586, fourFunc_wire_563_14);
notg #(0, 0) NOT_35 (fourFunc_wire_587, fourFunc_wire_563_15);
notg #(0, 0) NOT_36 (fourFunc_wire_588, fourFunc_wire_563_16);
notg #(0, 0) NOT_37 (fourFunc_wire_589, fourFunc_wire_563_17);
notg #(0, 0) NOT_38 (fourFunc_wire_590, fourFunc_wire_563_18);
notg #(0, 0) NOT_39 (fourFunc_wire_591, fourFunc_wire_563_19);
or_n #(2, 0, 0) OR_137 (fourFunc_wire_592, {fourFunc_wire_582, fourFunc_wire_593_0});
or_n #(2, 0, 0) OR_138 (fourFunc_wire_594, {fourFunc_wire_595, fourFunc_wire_593_1});
notg #(0, 0) NOT_40 (fourFunc_wire_596, fourFunc_wire_597);
and_n #(2, 0, 0) AND_226 (fourFunc_wire_595, {fourFunc_wire_596, fourFunc_wire_598_0});
or_n #(4, 0, 0) OR_139 (fourFunc_wire_599, {fourFunc_wire_600_0, fourFunc_wire_601_0, fourFunc_wire_602_0, fourFunc_wire_598_1});
and_n #(2, 0, 0) AND_227 (fourFunc_wire_439, {fourFunc_wire_11_10, fourFunc_wire_2_16});
and_n #(3, 0, 0) AND_228 (fourFunc_wire_612, {fourFunc_wire_11_11, fourFunc_wire_2_17, fourFunc_wire_3_12});
notg #(0, 0) NOT_41 (fourFunc_wire_613, fourFunc_wire_11_12);
and_n #(2, 0, 0) AND_229 (fourFunc_wire_614, {fourFunc_wire_615, fourFunc_wire_616});
or_n #(2, 0, 0) OR_140 (fourFunc_wire_616, {fourFunc_wire_613, fourFunc_wire_617_0});
notg #(0, 0) NOT_42 (fourFunc_wire_615, fourFunc_wire_611_0);
or_n #(3, 0, 0) OR_141 (fourFunc_wire_618, {fourFunc_wire_617_1, fourFunc_wire_601_1, fourFunc_wire_611_1});
and_n #(2, 0, 0) AND_230 (fourFunc_wire_619, {fourFunc_wire_620, fourFunc_wire_440});
notg #(0, 0) NOT_43 (fourFunc_wire_620, fourFunc_wire_621_0);
or_n #(2, 0, 0) OR_142 (fourFunc_wire_622, {fourFunc_wire_621_1, fourFunc_wire_601_2});
and_n #(2, 0, 0) AND_231 (fourFunc_wire_623, {fourFunc_wire_624, fourFunc_wire_438});
notg #(0, 0) NOT_44 (fourFunc_wire_624, fourFunc_wire_621_2);
or_n #(2, 0, 0) OR_143 (fourFunc_wire_621, {fourFunc_wire_617_2, fourFunc_wire_611_2});
and_n #(2, 0, 0) AND_232 (fourFunc_wire_625, {fourFunc_wire_7_15, fourFunc_wire_617_3});
notg #(0, 0) NOT_45 (fourFunc_wire_626, fourFunc_wire_7_16);
notg #(0, 0) NOT_46 (fourFunc_wire_627, fourFunc_wire_7_17);
notg #(0, 0) NOT_47 (fourFunc_wire_628, fourFunc_wire_7_18);
notg #(0, 0) NOT_48 (fourFunc_wire_629, fourFunc_wire_7_19);
notg #(0, 0) NOT_49 (fourFunc_wire_630, fourFunc_wire_7_20);
notg #(0, 0) NOT_50 (fourFunc_wire_631, fourFunc_wire_7_21);
notg #(0, 0) NOT_51 (fourFunc_wire_632, fourFunc_wire_7_22);
notg #(0, 0) NOT_52 (fourFunc_wire_633, fourFunc_wire_7_23);
or_n #(2, 0, 0) OR_144 (fourFunc_wire_634, {fourFunc_wire_7_24, fourFunc_wire_635_0});
or_n #(2, 0, 0) OR_145 (fourFunc_wire_636, {fourFunc_wire_7_25, fourFunc_wire_637_0});
or_n #(2, 0, 0) OR_146 (fourFunc_wire_638, {fourFunc_wire_7_26, fourFunc_wire_639_0});
or_n #(2, 0, 0) OR_147 (fourFunc_wire_640, {fourFunc_wire_7_27, fourFunc_wire_641_0});
or_n #(2, 0, 0) OR_148 (fourFunc_wire_642, {fourFunc_wire_7_28, fourFunc_wire_643_0});
or_n #(2, 0, 0) OR_149 (fourFunc_wire_644, {fourFunc_wire_7_29, fourFunc_wire_645_0});
or_n #(2, 0, 0) OR_150 (fourFunc_wire_646, {fourFunc_wire_7_30, fourFunc_wire_647_0});
or_n #(2, 0, 0) OR_151 (fourFunc_wire_648, {fourFunc_wire_7_31, fourFunc_wire_649_0});
and_n #(2, 0, 0) AND_233 (fourFunc_wire_617, {fourFunc_wire_593_2, fourFunc_wire_650_0});
notg #(0, 0) NOT_53 (fourFunc_wire_651, fourFunc_wire_617_4);
notg #(0, 0) NOT_54 (fourFunc_wire_652, fourFunc_wire_617_5);
notg #(0, 0) NOT_55 (fourFunc_wire_653, fourFunc_wire_617_6);
and_n #(2, 0, 0) AND_234 (fourFunc_wire_654, {fourFunc_wire_617_7, fourFunc_wire_637_1});
notg #(0, 0) NOT_56 (fourFunc_wire_655, fourFunc_wire_617_8);
and_n #(2, 0, 0) AND_235 (fourFunc_wire_656, {fourFunc_wire_617_9, fourFunc_wire_641_1});
notg #(0, 0) NOT_57 (fourFunc_wire_657, fourFunc_wire_617_10);
and_n #(2, 0, 0) AND_236 (fourFunc_wire_658, {fourFunc_wire_617_11, fourFunc_wire_635_1});
or_n #(3, 0, 0) OR_152 (fourFunc_wire_659, {fourFunc_wire_617_12, fourFunc_wire_600_1, fourFunc_wire_611_3});
notg #(0, 0) NOT_58 (fourFunc_wire_660, fourFunc_wire_617_13);
and_n #(2, 0, 0) AND_237 (fourFunc_wire_661, {fourFunc_wire_617_14, fourFunc_wire_639_1});
notg #(0, 0) NOT_59 (fourFunc_wire_662, fourFunc_wire_617_15);
and_n #(2, 0, 0) AND_238 (fourFunc_wire_663, {fourFunc_wire_617_16, fourFunc_wire_643_1});
notg #(0, 0) NOT_60 (fourFunc_wire_664, fourFunc_wire_617_17);
and_n #(2, 0, 0) AND_239 (fourFunc_wire_665, {fourFunc_wire_617_18, fourFunc_wire_649_1});
notg #(0, 0) NOT_61 (fourFunc_wire_666, fourFunc_wire_617_19);
and_n #(2, 0, 0) AND_240 (fourFunc_wire_667, {fourFunc_wire_617_20, fourFunc_wire_645_1});
notg #(0, 0) NOT_62 (fourFunc_wire_668, fourFunc_wire_617_21);
and_n #(2, 0, 0) AND_241 (fourFunc_wire_669, {fourFunc_wire_617_22, fourFunc_wire_647_1});
notg #(0, 0) NOT_63 (fourFunc_wire_670, fourFunc_wire_617_23);
and_n #(2, 0, 0) AND_242 (fourFunc_wire_671, {fourFunc_wire_617_24, fourFunc_wire_634});
notg #(0, 0) NOT_64 (fourFunc_wire_672, fourFunc_wire_617_25);
and_n #(2, 0, 0) AND_243 (fourFunc_wire_673, {fourFunc_wire_617_26, fourFunc_wire_636});
notg #(0, 0) NOT_65 (fourFunc_wire_674, fourFunc_wire_617_27);
and_n #(2, 0, 0) AND_244 (fourFunc_wire_675, {fourFunc_wire_617_28, fourFunc_wire_638});
notg #(0, 0) NOT_66 (fourFunc_wire_676, fourFunc_wire_617_29);
and_n #(2, 0, 0) AND_245 (fourFunc_wire_677, {fourFunc_wire_617_30, fourFunc_wire_640});
notg #(0, 0) NOT_67 (fourFunc_wire_678, fourFunc_wire_617_31);
and_n #(2, 0, 0) AND_246 (fourFunc_wire_679, {fourFunc_wire_617_32, fourFunc_wire_642});
notg #(0, 0) NOT_68 (fourFunc_wire_680, fourFunc_wire_617_33);
and_n #(2, 0, 0) AND_247 (fourFunc_wire_681, {fourFunc_wire_617_34, fourFunc_wire_644});
notg #(0, 0) NOT_69 (fourFunc_wire_682, fourFunc_wire_617_35);
and_n #(2, 0, 0) AND_248 (fourFunc_wire_683, {fourFunc_wire_617_36, fourFunc_wire_646});
notg #(0, 0) NOT_70 (fourFunc_wire_684, fourFunc_wire_617_37);
and_n #(2, 0, 0) AND_249 (fourFunc_wire_685, {fourFunc_wire_617_38, fourFunc_wire_648});
or_n #(2, 0, 0) OR_153 (fourFunc_wire_431, {fourFunc_wire_686, fourFunc_wire_687});
and_n #(2, 0, 0) AND_250 (fourFunc_wire_686, {fourFunc_wire_598_2, fourFunc_wire_4});
notg #(0, 0) NOT_71 (fourFunc_wire_688, fourFunc_wire_598_3);
and_n #(2, 0, 0) AND_251 (fourFunc_wire_687, {fourFunc_wire_688, fourFunc_wire_564_0});
or_n #(2, 0, 0) OR_154 (fourFunc_wire_429, {fourFunc_wire_689, fourFunc_wire_690});
and_n #(2, 0, 0) AND_252 (fourFunc_wire_689, {fourFunc_wire_598_4, fourFunc_wire_17});
notg #(0, 0) NOT_72 (fourFunc_wire_691, fourFunc_wire_598_5);
and_n #(2, 0, 0) AND_253 (fourFunc_wire_690, {fourFunc_wire_691, fourFunc_wire_565_0});
or_n #(2, 0, 0) OR_155 (fourFunc_wire_428, {fourFunc_wire_692, fourFunc_wire_693});
and_n #(2, 0, 0) AND_254 (fourFunc_wire_692, {fourFunc_wire_598_6, fourFunc_wire_27});
notg #(0, 0) NOT_73 (fourFunc_wire_694, fourFunc_wire_598_7);
and_n #(2, 0, 0) AND_255 (fourFunc_wire_693, {fourFunc_wire_694, fourFunc_wire_566_0});
or_n #(2, 0, 0) OR_156 (fourFunc_wire_427, {fourFunc_wire_695, fourFunc_wire_696});
and_n #(2, 0, 0) AND_256 (fourFunc_wire_695, {fourFunc_wire_598_8, fourFunc_wire_39});
notg #(0, 0) NOT_74 (fourFunc_wire_697, fourFunc_wire_598_9);
and_n #(2, 0, 0) AND_257 (fourFunc_wire_696, {fourFunc_wire_697, fourFunc_wire_567_0});
or_n #(2, 0, 0) OR_157 (fourFunc_wire_426, {fourFunc_wire_698, fourFunc_wire_699});
and_n #(2, 0, 0) AND_258 (fourFunc_wire_698, {fourFunc_wire_598_10, fourFunc_wire_44});
notg #(0, 0) NOT_75 (fourFunc_wire_700, fourFunc_wire_598_11);
and_n #(2, 0, 0) AND_259 (fourFunc_wire_699, {fourFunc_wire_700, fourFunc_wire_568_0});
or_n #(2, 0, 0) OR_158 (fourFunc_wire_425, {fourFunc_wire_701, fourFunc_wire_702});
and_n #(2, 0, 0) AND_260 (fourFunc_wire_701, {fourFunc_wire_598_12, fourFunc_wire_46});
notg #(0, 0) NOT_76 (fourFunc_wire_703, fourFunc_wire_598_13);
and_n #(2, 0, 0) AND_261 (fourFunc_wire_702, {fourFunc_wire_703, fourFunc_wire_569_0});
or_n #(2, 0, 0) OR_159 (fourFunc_wire_424, {fourFunc_wire_704, fourFunc_wire_705});
and_n #(2, 0, 0) AND_262 (fourFunc_wire_704, {fourFunc_wire_598_14, fourFunc_wire_53});
notg #(0, 0) NOT_77 (fourFunc_wire_706, fourFunc_wire_598_15);
and_n #(2, 0, 0) AND_263 (fourFunc_wire_705, {fourFunc_wire_706, fourFunc_wire_570_0});
or_n #(2, 0, 0) OR_160 (fourFunc_wire_423, {fourFunc_wire_707, fourFunc_wire_708});
and_n #(2, 0, 0) AND_264 (fourFunc_wire_707, {fourFunc_wire_598_16, fourFunc_wire_51});
notg #(0, 0) NOT_78 (fourFunc_wire_709, fourFunc_wire_598_17);
and_n #(2, 0, 0) AND_265 (fourFunc_wire_708, {fourFunc_wire_709, fourFunc_wire_571_0});
and_n #(2, 0, 0) AND_266 (fourFunc_wire_710, {fourFunc_wire_249, fourFunc_wire_676});
and_n #(2, 0, 0) AND_267 (fourFunc_wire_711, {fourFunc_wire_245, fourFunc_wire_670});
and_n #(2, 0, 0) AND_268 (fourFunc_wire_712, {fourFunc_wire_241, fourFunc_wire_678});
and_n #(2, 0, 0) AND_269 (fourFunc_wire_713, {fourFunc_wire_237, fourFunc_wire_680});
and_n #(2, 0, 0) AND_270 (fourFunc_wire_714, {fourFunc_wire_232, fourFunc_wire_682});
and_n #(2, 0, 0) AND_271 (fourFunc_wire_715, {fourFunc_wire_419, fourFunc_wire_684});
and_n #(2, 0, 0) AND_272 (fourFunc_wire_716, {fourFunc_wire_257, fourFunc_wire_672});
and_n #(2, 0, 0) AND_273 (fourFunc_wire_717, {fourFunc_wire_253, fourFunc_wire_674});
or_n #(2, 0, 0) OR_161 (fourFunc_wire_718, {fourFunc_wire_604, fourFunc_wire_611_4});
and_n #(2, 0, 0) AND_274 (fourFunc_wire_719, {fourFunc_wire_600_2, fourFunc_wire_612_0});
and_n #(2, 0, 0) AND_275 (fourFunc_wire_603, {fourFunc_wire_719, fourFunc_wire_720});
notg #(0, 0) NOT_79 (fourFunc_wire_720, fourFunc_wire_610_0);
and_n #(2, 0, 0) AND_276 (fourFunc_wire_721, {fourFunc_wire_600_3, fourFunc_wire_722});
notg #(0, 0) NOT_80 (fourFunc_wire_723, fourFunc_wire_610_1);
and_n #(2, 0, 0) AND_277 (fourFunc_wire_605, {fourFunc_wire_723, fourFunc_wire_601_3});
notg #(0, 0) NOT_81 (fourFunc_wire_724, fourFunc_wire_610_2);
and_n #(2, 0, 0) AND_278 (fourFunc_wire_606, {fourFunc_wire_724, fourFunc_wire_602_1});
notg #(0, 0) NOT_82 (fourFunc_wire_725, fourFunc_wire_610_3);
and_n #(2, 0, 0) AND_279 (fourFunc_wire_607, {fourFunc_wire_725, fourFunc_wire_598_18});
and_n #(2, 0, 0) AND_280 (fourFunc_wire_726, {fourFunc_wire_593_3, fourFunc_wire_650_1});
or_n #(2, 0, 0) OR_162 (fourFunc_wire_727, {fourFunc_wire_726, fourFunc_wire_721});
notg #(0, 0) NOT_83 (fourFunc_wire_722, fourFunc_wire_612_1);
notg #(0, 0) NOT_84 (fourFunc_wire_728, fourFunc_wire_610_4);
and_n #(2, 0, 0) AND_281 (fourFunc_wire_608, {fourFunc_wire_728, fourFunc_wire_727});
and_n #(2, 0, 0) AND_282 (fourFunc_wire_729, {fourFunc_wire_593_4, fourFunc_wire_730});
or_n #(2, 0, 0) OR_163 (fourFunc_wire_731, {fourFunc_wire_718, fourFunc_wire_729});
notg #(0, 0) NOT_85 (fourFunc_wire_730, fourFunc_wire_650_2);
notg #(0, 0) NOT_86 (fourFunc_wire_732, fourFunc_wire_610_5);
and_n #(2, 0, 0) AND_283 (fourFunc_wire_609, {fourFunc_wire_732, fourFunc_wire_731});
or_n #(2, 0, 0) OR_164 (fourFunc_wire_733, {fourFunc_wire_611_5, fourFunc_wire_734});
notg #(0, 0) NOT_87 (fourFunc_wire_735, fourFunc_wire_611_6);
notg #(0, 0) NOT_88 (fourFunc_wire_736, fourFunc_wire_611_7);
notg #(0, 0) NOT_89 (fourFunc_wire_737, fourFunc_wire_611_8);
notg #(0, 0) NOT_90 (fourFunc_wire_738, fourFunc_wire_611_9);
notg #(0, 0) NOT_91 (fourFunc_wire_739, fourFunc_wire_611_10);
notg #(0, 0) NOT_92 (fourFunc_wire_740, fourFunc_wire_611_11);
notg #(0, 0) NOT_93 (fourFunc_wire_741, fourFunc_wire_611_12);
notg #(0, 0) NOT_94 (fourFunc_wire_742, fourFunc_wire_611_13);
notg #(0, 0) NOT_95 (fourFunc_wire_743, fourFunc_wire_611_14);
notg #(0, 0) NOT_96 (fourFunc_wire_744, fourFunc_wire_611_15);
notg #(0, 0) NOT_97 (fourFunc_wire_745, fourFunc_wire_611_16);
notg #(0, 0) NOT_98 (fourFunc_wire_746, fourFunc_wire_611_17);
notg #(0, 0) NOT_99 (fourFunc_wire_747, fourFunc_wire_611_18);
notg #(0, 0) NOT_100 (fourFunc_wire_748, fourFunc_wire_611_19);
notg #(0, 0) NOT_101 (fourFunc_wire_749, fourFunc_wire_611_20);
notg #(0, 0) NOT_102 (fourFunc_wire_750, fourFunc_wire_611_21);
notg #(0, 0) NOT_103 (fourFunc_wire_751, fourFunc_wire_611_22);
notg #(0, 0) NOT_104 (fourFunc_wire_752, fourFunc_wire_611_23);
notg #(0, 0) NOT_105 (fourFunc_wire_753, fourFunc_wire_611_24);
notg #(0, 0) NOT_106 (fourFunc_wire_754, fourFunc_wire_611_25);
notg #(0, 0) NOT_107 (fourFunc_wire_755, fourFunc_wire_611_26);
notg #(0, 0) NOT_108 (fourFunc_wire_756, fourFunc_wire_611_27);
notg #(0, 0) NOT_109 (fourFunc_wire_757, fourFunc_wire_611_28);
notg #(0, 0) NOT_110 (fourFunc_wire_758, fourFunc_wire_611_29);
notg #(0, 0) NOT_111 (fourFunc_wire_759, fourFunc_wire_611_30);
notg #(0, 0) NOT_112 (fourFunc_wire_760, fourFunc_wire_611_31);
and_n #(2, 0, 0) AND_284 (fourFunc_wire_761, {fourFunc_wire_735, fourFunc_wire_637_2});
and_n #(2, 0, 0) AND_285 (fourFunc_wire_762, {fourFunc_wire_736, fourFunc_wire_639_2});
and_n #(2, 0, 0) AND_286 (fourFunc_wire_763, {fourFunc_wire_737, fourFunc_wire_641_2});
and_n #(2, 0, 0) AND_287 (fourFunc_wire_764, {fourFunc_wire_738, fourFunc_wire_635_2});
and_n #(2, 0, 0) AND_288 (fourFunc_wire_765, {fourFunc_wire_739, fourFunc_wire_643_2});
and_n #(2, 0, 0) AND_289 (fourFunc_wire_766, {fourFunc_wire_740, fourFunc_wire_645_2});
and_n #(2, 0, 0) AND_290 (fourFunc_wire_767, {fourFunc_wire_741, fourFunc_wire_647_2});
and_n #(2, 0, 0) AND_291 (fourFunc_wire_768, {fourFunc_wire_742, fourFunc_wire_649_2});
and_n #(2, 0, 0) AND_292 (fourFunc_wire_769, {fourFunc_wire_770, fourFunc_wire_745});
or_n #(2, 0, 0) OR_165 (fourFunc_wire_771, {fourFunc_wire_572, fourFunc_wire_772});
and_n #(2, 0, 0) AND_293 (fourFunc_wire_773, {fourFunc_wire_771, fourFunc_wire_653});
or_n #(2, 0, 0) OR_166 (fourFunc_wire_770, {fourFunc_wire_773, fourFunc_wire_774});
nor_n #(2, 0, 0) NOR_8 (fourFunc_wire_772, {fourFunc_wire_563_20, fourFunc_wire_441});
and_n #(2, 0, 0) AND_294 (fourFunc_wire_774, {fourFunc_wire_654, fourFunc_wire_626});
and_n #(2, 0, 0) AND_295 (fourFunc_wire_775, {fourFunc_wire_776, fourFunc_wire_748});
or_n #(2, 0, 0) OR_167 (fourFunc_wire_777, {fourFunc_wire_573, fourFunc_wire_778});
and_n #(2, 0, 0) AND_296 (fourFunc_wire_779, {fourFunc_wire_660, fourFunc_wire_777});
or_n #(2, 0, 0) OR_168 (fourFunc_wire_776, {fourFunc_wire_779, fourFunc_wire_780});
and_n #(2, 0, 0) AND_297 (fourFunc_wire_778, {fourFunc_wire_587, fourFunc_wire_473});
and_n #(2, 0, 0) AND_298 (fourFunc_wire_780, {fourFunc_wire_661, fourFunc_wire_629});
and_n #(2, 0, 0) AND_299 (fourFunc_wire_781, {fourFunc_wire_782, fourFunc_wire_746});
or_n #(2, 0, 0) OR_169 (fourFunc_wire_783, {fourFunc_wire_574, fourFunc_wire_784});
and_n #(2, 0, 0) AND_300 (fourFunc_wire_785, {fourFunc_wire_655, fourFunc_wire_783});
or_n #(2, 0, 0) OR_170 (fourFunc_wire_782, {fourFunc_wire_785, fourFunc_wire_786});
and_n #(2, 0, 0) AND_301 (fourFunc_wire_784, {fourFunc_wire_585, fourFunc_wire_469});
and_n #(2, 0, 0) AND_302 (fourFunc_wire_786, {fourFunc_wire_656, fourFunc_wire_627});
and_n #(2, 0, 0) AND_303 (fourFunc_wire_787, {fourFunc_wire_788, fourFunc_wire_747});
or_n #(2, 0, 0) OR_171 (fourFunc_wire_789, {fourFunc_wire_575, fourFunc_wire_790});
and_n #(2, 0, 0) AND_304 (fourFunc_wire_791, {fourFunc_wire_657, fourFunc_wire_789});
or_n #(2, 0, 0) OR_172 (fourFunc_wire_788, {fourFunc_wire_791, fourFunc_wire_792});
and_n #(2, 0, 0) AND_305 (fourFunc_wire_790, {fourFunc_wire_586, fourFunc_wire_465});
and_n #(2, 0, 0) AND_306 (fourFunc_wire_792, {fourFunc_wire_658, fourFunc_wire_628});
and_n #(2, 0, 0) AND_307 (fourFunc_wire_793, {fourFunc_wire_794, fourFunc_wire_749});
or_n #(2, 0, 0) OR_173 (fourFunc_wire_795, {fourFunc_wire_576, fourFunc_wire_796});
and_n #(2, 0, 0) AND_308 (fourFunc_wire_797, {fourFunc_wire_662, fourFunc_wire_795});
or_n #(2, 0, 0) OR_174 (fourFunc_wire_794, {fourFunc_wire_797, fourFunc_wire_798});
and_n #(2, 0, 0) AND_309 (fourFunc_wire_796, {fourFunc_wire_588, fourFunc_wire_461});
and_n #(2, 0, 0) AND_310 (fourFunc_wire_798, {fourFunc_wire_663, fourFunc_wire_630});
and_n #(2, 0, 0) AND_311 (fourFunc_wire_799, {fourFunc_wire_800, fourFunc_wire_751});
or_n #(2, 0, 0) OR_175 (fourFunc_wire_801, {fourFunc_wire_577, fourFunc_wire_802});
and_n #(2, 0, 0) AND_312 (fourFunc_wire_803, {fourFunc_wire_666, fourFunc_wire_801});
or_n #(2, 0, 0) OR_176 (fourFunc_wire_800, {fourFunc_wire_803, fourFunc_wire_804});
and_n #(2, 0, 0) AND_313 (fourFunc_wire_802, {fourFunc_wire_590, fourFunc_wire_457});
and_n #(2, 0, 0) AND_314 (fourFunc_wire_804, {fourFunc_wire_667, fourFunc_wire_632});
and_n #(2, 0, 0) AND_315 (fourFunc_wire_805, {fourFunc_wire_806, fourFunc_wire_752});
or_n #(2, 0, 0) OR_177 (fourFunc_wire_807, {fourFunc_wire_578, fourFunc_wire_808});
and_n #(2, 0, 0) AND_316 (fourFunc_wire_809, {fourFunc_wire_668, fourFunc_wire_807});
or_n #(2, 0, 0) OR_178 (fourFunc_wire_806, {fourFunc_wire_809, fourFunc_wire_810});
and_n #(2, 0, 0) AND_317 (fourFunc_wire_808, {fourFunc_wire_591, fourFunc_wire_453});
and_n #(2, 0, 0) AND_318 (fourFunc_wire_810, {fourFunc_wire_669, fourFunc_wire_633});
and_n #(2, 0, 0) AND_319 (fourFunc_wire_811, {fourFunc_wire_812, fourFunc_wire_750});
or_n #(2, 0, 0) OR_179 (fourFunc_wire_813, {fourFunc_wire_579, fourFunc_wire_814});
and_n #(2, 0, 0) AND_320 (fourFunc_wire_815, {fourFunc_wire_664, fourFunc_wire_813});
or_n #(2, 0, 0) OR_180 (fourFunc_wire_812, {fourFunc_wire_815, fourFunc_wire_816});
and_n #(2, 0, 0) AND_321 (fourFunc_wire_814, {fourFunc_wire_589, fourFunc_wire_449});
and_n #(2, 0, 0) AND_322 (fourFunc_wire_816, {fourFunc_wire_665, fourFunc_wire_631});
and_n #(2, 0, 0) AND_323 (fourFunc_wire_817, {fourFunc_wire_743, fourFunc_wire_818});
or_n #(2, 0, 0) OR_181 (fourFunc_wire_818, {fourFunc_wire_625, fourFunc_wire_819});
or_n #(2, 0, 0) OR_182 (fourFunc_wire_820, {fourFunc_wire_580, fourFunc_wire_821});
and_n #(2, 0, 0) AND_324 (fourFunc_wire_821, {fourFunc_wire_583, fourFunc_wire_446});
and_n #(2, 0, 0) AND_325 (fourFunc_wire_819, {fourFunc_wire_651, fourFunc_wire_820});
and_n #(3, 0, 0) AND_326 (fourFunc_wire_822, {fourFunc_wire_744, fourFunc_wire_652, fourFunc_wire_823});
or_n #(2, 0, 0) OR_183 (fourFunc_wire_823, {fourFunc_wire_581, fourFunc_wire_824});
and_n #(2, 0, 0) AND_327 (fourFunc_wire_824, {fourFunc_wire_584, fourFunc_wire_443});
and_n #(2, 0, 0) AND_328 (fourFunc_wire_825, {fourFunc_wire_754, fourFunc_wire_826});
or_n #(2, 0, 0) OR_184 (fourFunc_wire_826, {fourFunc_wire_673, fourFunc_wire_716});
notg #(0, 0) NOT_113 (fourFunc_wire_734, fourFunc_wire_827);
and_n #(2, 0, 0) AND_329 (fourFunc_wire_828, {fourFunc_wire_755, fourFunc_wire_829});
or_n #(2, 0, 0) OR_185 (fourFunc_wire_829, {fourFunc_wire_675, fourFunc_wire_717});
and_n #(2, 0, 0) AND_330 (fourFunc_wire_830, {fourFunc_wire_756, fourFunc_wire_831});
or_n #(2, 0, 0) OR_186 (fourFunc_wire_831, {fourFunc_wire_677, fourFunc_wire_710});
and_n #(2, 0, 0) AND_331 (fourFunc_wire_832, {fourFunc_wire_753, fourFunc_wire_833});
or_n #(2, 0, 0) OR_187 (fourFunc_wire_833, {fourFunc_wire_671, fourFunc_wire_711});
and_n #(2, 0, 0) AND_332 (fourFunc_wire_834, {fourFunc_wire_757, fourFunc_wire_835});
or_n #(2, 0, 0) OR_188 (fourFunc_wire_835, {fourFunc_wire_679, fourFunc_wire_712});
and_n #(2, 0, 0) AND_333 (fourFunc_wire_836, {fourFunc_wire_758, fourFunc_wire_837});
or_n #(2, 0, 0) OR_189 (fourFunc_wire_837, {fourFunc_wire_681, fourFunc_wire_713});
and_n #(2, 0, 0) AND_334 (fourFunc_wire_838, {fourFunc_wire_759, fourFunc_wire_839});
or_n #(2, 0, 0) OR_190 (fourFunc_wire_839, {fourFunc_wire_683, fourFunc_wire_714});
and_n #(2, 0, 0) AND_335 (fourFunc_wire_840, {fourFunc_wire_760, fourFunc_wire_841});
or_n #(2, 0, 0) OR_191 (fourFunc_wire_841, {fourFunc_wire_685, fourFunc_wire_715});
nor_n #(4, 0, 0) NOR_9 (fourFunc_wire_827, {fourFunc_wire_617_39, fourFunc_wire_602_2, fourFunc_wire_601_4, fourFunc_wire_598_19});
bufg #(0, 0) BUF_10 (busy_net_0, fourFunc_wire_599);
bufg #(0, 0) BUF_11 (fourFunc_wire_562, clk_net_0);
bufg #(0, 0) BUF_12 (fourFunc_wire_7, func_1);
bufg #(0, 0) BUF_13 (fourFunc_wire_597, func_0);
bufg #(0, 0) BUF_14 (resultFPart_7, fourFunc_wire_442_4);
bufg #(0, 0) BUF_15 (resultFPart_6, fourFunc_wire_476_6);
bufg #(0, 0) BUF_16 (resultFPart_5, fourFunc_wire_472_6);
bufg #(0, 0) BUF_17 (resultFPart_4, fourFunc_wire_468_6);
bufg #(0, 0) BUF_18 (resultFPart_3, fourFunc_wire_464_6);
bufg #(0, 0) BUF_19 (resultFPart_2, fourFunc_wire_460_6);
bufg #(0, 0) BUF_20 (resultFPart_1, fourFunc_wire_456_6);
bufg #(0, 0) BUF_21 (resultFPart_0, fourFunc_wire_452_6);
bufg #(0, 0) BUF_22 (resultIPart_1, fourFunc_wire_447_5);
bufg #(0, 0) BUF_23 (resultIPart_0, fourFunc_wire_444_2);
bufg #(0, 0) BUF_24 (fourFunc_wire_610, rst_net_0);
bufg #(0, 0) BUF_25 (fourFunc_wire_650, start_net_0);
bufg #(0, 0) BUF_26 (fourFunc_wire_637, x_7);
bufg #(0, 0) BUF_27 (fourFunc_wire_639, x_6);
bufg #(0, 0) BUF_28 (fourFunc_wire_641, x_5);
bufg #(0, 0) BUF_29 (fourFunc_wire_635, x_4);
bufg #(0, 0) BUF_30 (fourFunc_wire_643, x_3);
bufg #(0, 0) BUF_31 (fourFunc_wire_645, x_2);
bufg #(0, 0) BUF_32 (fourFunc_wire_647, x_1);
bufg #(0, 0) BUF_33 (fourFunc_wire_649, x_0);
and_n #(2, 0, 0) AND_336 (NOT_intermediateXXXwire_721_AND_intermediateXXXwire_718, {fourFunc_wire_563_21, NOT_intermediateXXXwire_721});
and_n #(2, 0, 0) AND_337 (fourFunc_wire_842, {fourFunc_wire_594_0, fourFunc_wire_592});
or_n #(2, 0, 0) OR_192 (NOT_intermediateXXXwire_721_AND_intermediateXXXwire_718_OR_intermediateXXXwire_721_AND_intermediateXXXwire_719, {NOT_intermediateXXXwire_721_AND_intermediateXXXwire_718, fourFunc_wire_842});
notg #(0, 0) NOT_114 (NOT_intermediateXXXwire_721, fourFunc_wire_594_1);
and_n #(2, 0, 0) AND_338 (NOT_intermediateXXXwire_731_AND_intermediateXXXwire_61, {fourFunc_wire_11_13, NOT_intermediateXXXwire_731});
and_n #(2, 0, 0) AND_339 (fourFunc_wire_843, {fourFunc_wire_618_0, fourFunc_wire_614});
or_n #(2, 0, 0) OR_193 (NOT_intermediateXXXwire_731_AND_intermediateXXXwire_61_OR_intermediateXXXwire_731_AND_intermediateXXXwire_727, {NOT_intermediateXXXwire_731_AND_intermediateXXXwire_61, fourFunc_wire_843});
notg #(0, 0) NOT_115 (NOT_intermediateXXXwire_731, fourFunc_wire_618_1);
and_n #(2, 0, 0) AND_340 (NOT_intermediateXXXwire_735_AND_intermediateXXXwire_63, {fourFunc_wire_3_13, NOT_intermediateXXXwire_735_0});
and_n #(2, 0, 0) AND_341 (fourFunc_wire_844, {fourFunc_wire_622_0, fourFunc_wire_623});
or_n #(2, 0, 0) OR_194 (NOT_intermediateXXXwire_735_AND_intermediateXXXwire_63_OR_intermediateXXXwire_735_AND_intermediateXXXwire_737, {NOT_intermediateXXXwire_735_AND_intermediateXXXwire_63, fourFunc_wire_844});
notg #(0, 0) NOT_116 (NOT_intermediateXXXwire_735, fourFunc_wire_622_1);
and_n #(2, 0, 0) AND_342 (NOT_intermediateXXXwire_735_AND_intermediateXXXwire_62, {fourFunc_wire_2_18, NOT_intermediateXXXwire_735_1});
and_n #(2, 0, 0) AND_343 (fourFunc_wire_845, {fourFunc_wire_622_2, fourFunc_wire_619});
or_n #(2, 0, 0) OR_195 (NOT_intermediateXXXwire_735_AND_intermediateXXXwire_62_OR_intermediateXXXwire_735_AND_intermediateXXXwire_733, {NOT_intermediateXXXwire_735_AND_intermediateXXXwire_62, fourFunc_wire_845});
and_n #(2, 0, 0) AND_344 (NOT_intermediateXXXwire_739_AND_intermediateXXXwire_796, {fourFunc_wire_564_1, NOT_intermediateXXXwire_739_0});
and_n #(2, 0, 0) AND_345 (fourFunc_wire_846, {fourFunc_wire_621_3, fourFunc_wire_761});
or_n #(2, 0, 0) OR_196 (NOT_intermediateXXXwire_739_AND_intermediateXXXwire_796_OR_intermediateXXXwire_739_AND_intermediateXXXwire_797, {NOT_intermediateXXXwire_739_AND_intermediateXXXwire_796, fourFunc_wire_846});
notg #(0, 0) NOT_117 (NOT_intermediateXXXwire_739, fourFunc_wire_621_4);
and_n #(2, 0, 0) AND_346 (NOT_intermediateXXXwire_739_AND_intermediateXXXwire_799, {fourFunc_wire_565_1, NOT_intermediateXXXwire_739_1});
and_n #(2, 0, 0) AND_347 (fourFunc_wire_847, {fourFunc_wire_621_5, fourFunc_wire_762});
or_n #(2, 0, 0) OR_197 (NOT_intermediateXXXwire_739_AND_intermediateXXXwire_799_OR_intermediateXXXwire_739_AND_intermediateXXXwire_800, {NOT_intermediateXXXwire_739_AND_intermediateXXXwire_799, fourFunc_wire_847});
and_n #(2, 0, 0) AND_348 (NOT_intermediateXXXwire_739_AND_intermediateXXXwire_802, {fourFunc_wire_566_1, NOT_intermediateXXXwire_739_2});
and_n #(2, 0, 0) AND_349 (fourFunc_wire_848, {fourFunc_wire_621_6, fourFunc_wire_763});
or_n #(2, 0, 0) OR_198 (NOT_intermediateXXXwire_739_AND_intermediateXXXwire_802_OR_intermediateXXXwire_739_AND_intermediateXXXwire_803, {NOT_intermediateXXXwire_739_AND_intermediateXXXwire_802, fourFunc_wire_848});
and_n #(2, 0, 0) AND_350 (NOT_intermediateXXXwire_739_AND_intermediateXXXwire_805, {fourFunc_wire_567_1, NOT_intermediateXXXwire_739_3});
and_n #(2, 0, 0) AND_351 (fourFunc_wire_849, {fourFunc_wire_621_7, fourFunc_wire_764});
or_n #(2, 0, 0) OR_199 (NOT_intermediateXXXwire_739_AND_intermediateXXXwire_805_OR_intermediateXXXwire_739_AND_intermediateXXXwire_806, {NOT_intermediateXXXwire_739_AND_intermediateXXXwire_805, fourFunc_wire_849});
and_n #(2, 0, 0) AND_352 (NOT_intermediateXXXwire_739_AND_intermediateXXXwire_808, {fourFunc_wire_568_1, NOT_intermediateXXXwire_739_4});
and_n #(2, 0, 0) AND_353 (fourFunc_wire_850, {fourFunc_wire_621_8, fourFunc_wire_765});
or_n #(2, 0, 0) OR_200 (NOT_intermediateXXXwire_739_AND_intermediateXXXwire_808_OR_intermediateXXXwire_739_AND_intermediateXXXwire_809, {NOT_intermediateXXXwire_739_AND_intermediateXXXwire_808, fourFunc_wire_850});
and_n #(2, 0, 0) AND_354 (NOT_intermediateXXXwire_739_AND_intermediateXXXwire_811, {fourFunc_wire_569_1, NOT_intermediateXXXwire_739_5});
and_n #(2, 0, 0) AND_355 (fourFunc_wire_851, {fourFunc_wire_621_9, fourFunc_wire_766});
or_n #(2, 0, 0) OR_201 (NOT_intermediateXXXwire_739_AND_intermediateXXXwire_811_OR_intermediateXXXwire_739_AND_intermediateXXXwire_812, {NOT_intermediateXXXwire_739_AND_intermediateXXXwire_811, fourFunc_wire_851});
and_n #(2, 0, 0) AND_356 (NOT_intermediateXXXwire_739_AND_intermediateXXXwire_814, {fourFunc_wire_570_1, NOT_intermediateXXXwire_739_6});
and_n #(2, 0, 0) AND_357 (fourFunc_wire_852, {fourFunc_wire_621_10, fourFunc_wire_767});
or_n #(2, 0, 0) OR_202 (NOT_intermediateXXXwire_739_AND_intermediateXXXwire_814_OR_intermediateXXXwire_739_AND_intermediateXXXwire_815, {NOT_intermediateXXXwire_739_AND_intermediateXXXwire_814, fourFunc_wire_852});
and_n #(2, 0, 0) AND_358 (NOT_intermediateXXXwire_739_AND_intermediateXXXwire_817, {fourFunc_wire_571_1, NOT_intermediateXXXwire_739_7});
and_n #(2, 0, 0) AND_359 (fourFunc_wire_853, {fourFunc_wire_621_11, fourFunc_wire_768});
or_n #(2, 0, 0) OR_203 (NOT_intermediateXXXwire_739_AND_intermediateXXXwire_817_OR_intermediateXXXwire_739_AND_intermediateXXXwire_818, {NOT_intermediateXXXwire_739_AND_intermediateXXXwire_817, fourFunc_wire_853});
and_n #(2, 0, 0) AND_360 (NOT_intermediateXXXwire_963_AND_intermediateXXXwire_955, {fourFunc_wire_422_11, NOT_intermediateXXXwire_963_0});
and_n #(2, 0, 0) AND_361 (fourFunc_wire_854, {fourFunc_wire_733_0, fourFunc_wire_825});
or_n #(2, 0, 0) OR_204 (NOT_intermediateXXXwire_963_AND_intermediateXXXwire_955_OR_intermediateXXXwire_963_AND_intermediateXXXwire_956, {NOT_intermediateXXXwire_963_AND_intermediateXXXwire_955, fourFunc_wire_854});
notg #(0, 0) NOT_118 (NOT_intermediateXXXwire_963, fourFunc_wire_733_1);
and_n #(2, 0, 0) AND_362 (NOT_intermediateXXXwire_963_AND_intermediateXXXwire_965, {fourFunc_wire_430_14, NOT_intermediateXXXwire_963_1});
and_n #(2, 0, 0) AND_363 (fourFunc_wire_855, {fourFunc_wire_733_2, fourFunc_wire_828});
or_n #(2, 0, 0) OR_205 (NOT_intermediateXXXwire_963_AND_intermediateXXXwire_965_OR_intermediateXXXwire_963_AND_intermediateXXXwire_966, {NOT_intermediateXXXwire_963_AND_intermediateXXXwire_965, fourFunc_wire_855});
and_n #(2, 0, 0) AND_364 (NOT_intermediateXXXwire_963_AND_intermediateXXXwire_973, {fourFunc_wire_432_14, NOT_intermediateXXXwire_963_2});
and_n #(2, 0, 0) AND_365 (fourFunc_wire_856, {fourFunc_wire_733_3, fourFunc_wire_830});
or_n #(2, 0, 0) OR_206 (NOT_intermediateXXXwire_963_AND_intermediateXXXwire_973_OR_intermediateXXXwire_963_AND_intermediateXXXwire_974, {NOT_intermediateXXXwire_963_AND_intermediateXXXwire_973, fourFunc_wire_856});
and_n #(2, 0, 0) AND_366 (NOT_intermediateXXXwire_963_AND_intermediateXXXwire_981, {fourFunc_wire_433_14, NOT_intermediateXXXwire_963_3});
and_n #(2, 0, 0) AND_367 (fourFunc_wire_857, {fourFunc_wire_733_4, fourFunc_wire_832});
or_n #(2, 0, 0) OR_207 (NOT_intermediateXXXwire_963_AND_intermediateXXXwire_981_OR_intermediateXXXwire_963_AND_intermediateXXXwire_982, {NOT_intermediateXXXwire_963_AND_intermediateXXXwire_981, fourFunc_wire_857});
and_n #(2, 0, 0) AND_368 (NOT_intermediateXXXwire_963_AND_intermediateXXXwire_989, {fourFunc_wire_434_14, NOT_intermediateXXXwire_963_4});
and_n #(2, 0, 0) AND_369 (fourFunc_wire_858, {fourFunc_wire_733_5, fourFunc_wire_834});
or_n #(2, 0, 0) OR_208 (NOT_intermediateXXXwire_963_AND_intermediateXXXwire_989_OR_intermediateXXXwire_963_AND_intermediateXXXwire_990, {NOT_intermediateXXXwire_963_AND_intermediateXXXwire_989, fourFunc_wire_858});
and_n #(2, 0, 0) AND_370 (NOT_intermediateXXXwire_963_AND_intermediateXXXwire_997, {fourFunc_wire_435_14, NOT_intermediateXXXwire_963_5});
and_n #(2, 0, 0) AND_371 (fourFunc_wire_859, {fourFunc_wire_733_6, fourFunc_wire_836});
or_n #(2, 0, 0) OR_209 (NOT_intermediateXXXwire_963_AND_intermediateXXXwire_997_OR_intermediateXXXwire_963_AND_intermediateXXXwire_998, {NOT_intermediateXXXwire_963_AND_intermediateXXXwire_997, fourFunc_wire_859});
and_n #(2, 0, 0) AND_372 (NOT_intermediateXXXwire_963_AND_intermediateXXXwire_1005, {fourFunc_wire_436_14, NOT_intermediateXXXwire_963_6});
and_n #(2, 0, 0) AND_373 (fourFunc_wire_860, {fourFunc_wire_733_7, fourFunc_wire_838});
or_n #(2, 0, 0) OR_210 (NOT_intermediateXXXwire_963_AND_intermediateXXXwire_1005_OR_intermediateXXXwire_963_AND_intermediateXXXwire_1006, {NOT_intermediateXXXwire_963_AND_intermediateXXXwire_1005, fourFunc_wire_860});
and_n #(2, 0, 0) AND_374 (NOT_intermediateXXXwire_963_AND_intermediateXXXwire_1013, {fourFunc_wire_437_14, NOT_intermediateXXXwire_963_7});
and_n #(2, 0, 0) AND_375 (fourFunc_wire_861, {fourFunc_wire_733_8, fourFunc_wire_840});
or_n #(2, 0, 0) OR_211 (NOT_intermediateXXXwire_963_AND_intermediateXXXwire_1013_OR_intermediateXXXwire_963_AND_intermediateXXXwire_1014, {NOT_intermediateXXXwire_963_AND_intermediateXXXwire_1013, fourFunc_wire_861});
and_n #(2, 0, 0) AND_376 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_820, {fourFunc_wire_442_5, NOT_intermediateXXXwire_834_0});
and_n #(2, 0, 0) AND_377 (fourFunc_wire_862, {fourFunc_wire_659_0, fourFunc_wire_769});
or_n #(2, 0, 0) OR_212 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_820_OR_intermediateXXXwire_834_AND_intermediateXXXwire_821, {NOT_intermediateXXXwire_834_AND_intermediateXXXwire_820, fourFunc_wire_862});
notg #(0, 0) NOT_119 (NOT_intermediateXXXwire_834, fourFunc_wire_659_1);
and_n #(2, 0, 0) AND_378 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_835, {fourFunc_wire_476_7, NOT_intermediateXXXwire_834_1});
and_n #(2, 0, 0) AND_379 (fourFunc_wire_863, {fourFunc_wire_659_2, fourFunc_wire_775});
or_n #(2, 0, 0) OR_213 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_835_OR_intermediateXXXwire_834_AND_intermediateXXXwire_836, {NOT_intermediateXXXwire_834_AND_intermediateXXXwire_835, fourFunc_wire_863});
and_n #(2, 0, 0) AND_380 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_848, {fourFunc_wire_472_7, NOT_intermediateXXXwire_834_2});
and_n #(2, 0, 0) AND_381 (fourFunc_wire_864, {fourFunc_wire_659_3, fourFunc_wire_781});
or_n #(2, 0, 0) OR_214 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_848_OR_intermediateXXXwire_834_AND_intermediateXXXwire_849, {NOT_intermediateXXXwire_834_AND_intermediateXXXwire_848, fourFunc_wire_864});
and_n #(2, 0, 0) AND_382 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_861, {fourFunc_wire_468_7, NOT_intermediateXXXwire_834_3});
and_n #(2, 0, 0) AND_383 (fourFunc_wire_865, {fourFunc_wire_659_4, fourFunc_wire_787});
or_n #(2, 0, 0) OR_215 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_861_OR_intermediateXXXwire_834_AND_intermediateXXXwire_862, {NOT_intermediateXXXwire_834_AND_intermediateXXXwire_861, fourFunc_wire_865});
and_n #(2, 0, 0) AND_384 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_874, {fourFunc_wire_464_7, NOT_intermediateXXXwire_834_4});
and_n #(2, 0, 0) AND_385 (fourFunc_wire_866, {fourFunc_wire_659_5, fourFunc_wire_793});
or_n #(2, 0, 0) OR_216 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_874_OR_intermediateXXXwire_834_AND_intermediateXXXwire_875, {NOT_intermediateXXXwire_834_AND_intermediateXXXwire_874, fourFunc_wire_866});
and_n #(2, 0, 0) AND_386 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_887, {fourFunc_wire_460_7, NOT_intermediateXXXwire_834_5});
and_n #(2, 0, 0) AND_387 (fourFunc_wire_867, {fourFunc_wire_659_6, fourFunc_wire_799});
or_n #(2, 0, 0) OR_217 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_887_OR_intermediateXXXwire_834_AND_intermediateXXXwire_888, {NOT_intermediateXXXwire_834_AND_intermediateXXXwire_887, fourFunc_wire_867});
and_n #(2, 0, 0) AND_388 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_900, {fourFunc_wire_456_7, NOT_intermediateXXXwire_834_6});
and_n #(2, 0, 0) AND_389 (fourFunc_wire_868, {fourFunc_wire_659_7, fourFunc_wire_805});
or_n #(2, 0, 0) OR_218 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_900_OR_intermediateXXXwire_834_AND_intermediateXXXwire_901, {NOT_intermediateXXXwire_834_AND_intermediateXXXwire_900, fourFunc_wire_868});
and_n #(2, 0, 0) AND_390 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_913, {fourFunc_wire_452_7, NOT_intermediateXXXwire_834_7});
and_n #(2, 0, 0) AND_391 (fourFunc_wire_869, {fourFunc_wire_659_8, fourFunc_wire_811});
or_n #(2, 0, 0) OR_219 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_913_OR_intermediateXXXwire_834_AND_intermediateXXXwire_914, {NOT_intermediateXXXwire_834_AND_intermediateXXXwire_913, fourFunc_wire_869});
and_n #(2, 0, 0) AND_392 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_926, {fourFunc_wire_447_6, NOT_intermediateXXXwire_834_8});
and_n #(2, 0, 0) AND_393 (fourFunc_wire_870, {fourFunc_wire_659_9, fourFunc_wire_817});
or_n #(2, 0, 0) OR_220 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_926_OR_intermediateXXXwire_834_AND_intermediateXXXwire_927, {NOT_intermediateXXXwire_834_AND_intermediateXXXwire_926, fourFunc_wire_870});
and_n #(2, 0, 0) AND_394 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_937, {fourFunc_wire_444_3, NOT_intermediateXXXwire_834_9});
and_n #(2, 0, 0) AND_395 (fourFunc_wire_871, {fourFunc_wire_659_10, fourFunc_wire_822});
or_n #(2, 0, 0) OR_221 (NOT_intermediateXXXwire_834_AND_intermediateXXXwire_937_OR_intermediateXXXwire_834_AND_intermediateXXXwire_938, {NOT_intermediateXXXwire_834_AND_intermediateXXXwire_937, fourFunc_wire_871});
/* dff DFF_1  (fourFunc_wire_563, NOT_intermediateXXXwire_721_AND_intermediateXXXwire_718_OR_intermediateXXXwire_721_AND_intermediateXXXwire_719, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_2  (fourFunc_wire_11, NOT_intermediateXXXwire_731_AND_intermediateXXXwire_61_OR_intermediateXXXwire_731_AND_intermediateXXXwire_727, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_3  (fourFunc_wire_3, NOT_intermediateXXXwire_735_AND_intermediateXXXwire_63_OR_intermediateXXXwire_735_AND_intermediateXXXwire_737, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_4  (fourFunc_wire_2, NOT_intermediateXXXwire_735_AND_intermediateXXXwire_62_OR_intermediateXXXwire_735_AND_intermediateXXXwire_733, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_5  (fourFunc_wire_564, NOT_intermediateXXXwire_739_AND_intermediateXXXwire_796_OR_intermediateXXXwire_739_AND_intermediateXXXwire_797, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_6  (fourFunc_wire_565, NOT_intermediateXXXwire_739_AND_intermediateXXXwire_799_OR_intermediateXXXwire_739_AND_intermediateXXXwire_800, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_7  (fourFunc_wire_566, NOT_intermediateXXXwire_739_AND_intermediateXXXwire_802_OR_intermediateXXXwire_739_AND_intermediateXXXwire_803, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_8  (fourFunc_wire_567, NOT_intermediateXXXwire_739_AND_intermediateXXXwire_805_OR_intermediateXXXwire_739_AND_intermediateXXXwire_806, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_9  (fourFunc_wire_568, NOT_intermediateXXXwire_739_AND_intermediateXXXwire_808_OR_intermediateXXXwire_739_AND_intermediateXXXwire_809, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_10  (fourFunc_wire_569, NOT_intermediateXXXwire_739_AND_intermediateXXXwire_811_OR_intermediateXXXwire_739_AND_intermediateXXXwire_812, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_11  (fourFunc_wire_570, NOT_intermediateXXXwire_739_AND_intermediateXXXwire_814_OR_intermediateXXXwire_739_AND_intermediateXXXwire_815, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_12  (fourFunc_wire_571, NOT_intermediateXXXwire_739_AND_intermediateXXXwire_817_OR_intermediateXXXwire_739_AND_intermediateXXXwire_818, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_13  (fourFunc_wire_422, NOT_intermediateXXXwire_963_AND_intermediateXXXwire_955_OR_intermediateXXXwire_963_AND_intermediateXXXwire_956, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_14  (fourFunc_wire_430, NOT_intermediateXXXwire_963_AND_intermediateXXXwire_965_OR_intermediateXXXwire_963_AND_intermediateXXXwire_966, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_15  (fourFunc_wire_432, NOT_intermediateXXXwire_963_AND_intermediateXXXwire_973_OR_intermediateXXXwire_963_AND_intermediateXXXwire_974, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_16  (fourFunc_wire_433, NOT_intermediateXXXwire_963_AND_intermediateXXXwire_981_OR_intermediateXXXwire_963_AND_intermediateXXXwire_982, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_17  (fourFunc_wire_434, NOT_intermediateXXXwire_963_AND_intermediateXXXwire_989_OR_intermediateXXXwire_963_AND_intermediateXXXwire_990, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_18  (fourFunc_wire_435, NOT_intermediateXXXwire_963_AND_intermediateXXXwire_997_OR_intermediateXXXwire_963_AND_intermediateXXXwire_998, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_19  (fourFunc_wire_436, NOT_intermediateXXXwire_963_AND_intermediateXXXwire_1005_OR_intermediateXXXwire_963_AND_intermediateXXXwire_1006, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_20  (fourFunc_wire_437, NOT_intermediateXXXwire_963_AND_intermediateXXXwire_1013_OR_intermediateXXXwire_963_AND_intermediateXXXwire_1014, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_21  (fourFunc_wire_442, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_820_OR_intermediateXXXwire_834_AND_intermediateXXXwire_821, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_22  (fourFunc_wire_476, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_835_OR_intermediateXXXwire_834_AND_intermediateXXXwire_836, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_23  (fourFunc_wire_472, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_848_OR_intermediateXXXwire_834_AND_intermediateXXXwire_849, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_24  (fourFunc_wire_468, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_861_OR_intermediateXXXwire_834_AND_intermediateXXXwire_862, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_25  (fourFunc_wire_464, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_874_OR_intermediateXXXwire_834_AND_intermediateXXXwire_875, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_26  (fourFunc_wire_460, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_887_OR_intermediateXXXwire_834_AND_intermediateXXXwire_888, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_27  (fourFunc_wire_456, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_900_OR_intermediateXXXwire_834_AND_intermediateXXXwire_901, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_28  (fourFunc_wire_452, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_913_OR_intermediateXXXwire_834_AND_intermediateXXXwire_914, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_29  (fourFunc_wire_447, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_926_OR_intermediateXXXwire_834_AND_intermediateXXXwire_927, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_30  (fourFunc_wire_444, NOT_intermediateXXXwire_834_AND_intermediateXXXwire_937_OR_intermediateXXXwire_834_AND_intermediateXXXwire_938, fourFunc_wire_562, fourFunc_wire_561, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_31  (fourFunc_wire_604, fourFunc_wire_603, fourFunc_wire_562, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_32  (fourFunc_wire_600, fourFunc_wire_605, fourFunc_wire_562, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_33  (fourFunc_wire_601, fourFunc_wire_606, fourFunc_wire_562, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_34  (fourFunc_wire_602, fourFunc_wire_607, fourFunc_wire_562, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_35  (fourFunc_wire_598, fourFunc_wire_608, fourFunc_wire_562, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_36  (fourFunc_wire_593, fourFunc_wire_609, fourFunc_wire_562, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_37  (fourFunc_wire_611, fourFunc_wire_610, fourFunc_wire_562, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
 */
endmodule
